
module Cipher ( clk, rst, EncDec, Input, Key, Tweak, Output, done );
  input [63:0] Input;
  input [127:0] Key;
  input [63:0] Tweak;
  output [63:0] Output;
  input clk, rst, EncDec;
  output done;
  wire   selectsReg_0_, selectsNext_0_, n3, n4, n5, n6, n7,
         MCInst_XOR_r0_Inst_0_n5, MCInst_XOR_r0_Inst_1_n5,
         MCInst_XOR_r0_Inst_2_n5, MCInst_XOR_r0_Inst_3_n5,
         MCInst_XOR_r0_Inst_4_n5, MCInst_XOR_r0_Inst_5_n5,
         MCInst_XOR_r0_Inst_6_n5, MCInst_XOR_r0_Inst_7_n5,
         MCInst_XOR_r0_Inst_8_n5, MCInst_XOR_r0_Inst_9_n5,
         MCInst_XOR_r0_Inst_10_n5, MCInst_XOR_r0_Inst_11_n5,
         MCInst_XOR_r0_Inst_12_n5, MCInst_XOR_r0_Inst_13_n5,
         MCInst_XOR_r0_Inst_14_n5, MCInst_XOR_r0_Inst_15_n5,
         AddKeyConstXOR_XORInst_0_0_n5, AddKeyConstXOR_XORInst_0_1_n5,
         AddKeyConstXOR_XORInst_0_2_n5, AddKeyConstXOR_XORInst_1_0_n5,
         AddKeyConstXOR_XORInst_1_1_n5, AddKeyConstXOR_XORInst_1_2_n5,
         AddKeyConstXOR_XORInst_1_3_n5,
         F_StateRegOutput_Inst_LFInst_0_LFInst_0_n3,
         F_StateRegOutput_Inst_LFInst_0_LFInst_1_n3,
         F_StateRegOutput_Inst_LFInst_1_LFInst_0_n3,
         F_StateRegOutput_Inst_LFInst_1_LFInst_1_n3,
         F_StateRegOutput_Inst_LFInst_2_LFInst_0_n3,
         F_StateRegOutput_Inst_LFInst_2_LFInst_1_n3,
         F_StateRegOutput_Inst_LFInst_3_LFInst_0_n3,
         F_StateRegOutput_Inst_LFInst_3_LFInst_1_n3,
         F_StateRegOutput_Inst_LFInst_4_LFInst_0_n3,
         F_StateRegOutput_Inst_LFInst_4_LFInst_1_n3,
         F_StateRegOutput_Inst_LFInst_5_LFInst_0_n3,
         F_StateRegOutput_Inst_LFInst_5_LFInst_1_n3,
         F_StateRegOutput_Inst_LFInst_6_LFInst_0_n3,
         F_StateRegOutput_Inst_LFInst_6_LFInst_1_n3,
         F_StateRegOutput_Inst_LFInst_7_LFInst_0_n3,
         F_StateRegOutput_Inst_LFInst_7_LFInst_1_n3,
         F_StateRegOutput_Inst_LFInst_8_LFInst_0_n3,
         F_StateRegOutput_Inst_LFInst_8_LFInst_1_n3,
         F_StateRegOutput_Inst_LFInst_9_LFInst_0_n3,
         F_StateRegOutput_Inst_LFInst_9_LFInst_1_n3,
         F_StateRegOutput_Inst_LFInst_10_LFInst_0_n3,
         F_StateRegOutput_Inst_LFInst_10_LFInst_1_n3,
         F_StateRegOutput_Inst_LFInst_11_LFInst_0_n3,
         F_StateRegOutput_Inst_LFInst_11_LFInst_1_n3,
         F_StateRegOutput_Inst_LFInst_12_LFInst_0_n3,
         F_StateRegOutput_Inst_LFInst_12_LFInst_1_n3,
         F_StateRegOutput_Inst_LFInst_13_LFInst_0_n3,
         F_StateRegOutput_Inst_LFInst_13_LFInst_1_n3,
         F_StateRegOutput_Inst_LFInst_14_LFInst_0_n3,
         F_StateRegOutput_Inst_LFInst_14_LFInst_1_n3,
         F_StateRegOutput_Inst_LFInst_15_LFInst_0_n3,
         F_StateRegOutput_Inst_LFInst_15_LFInst_1_n3,
         CipherErrorVecGen_XORInst_0_3_n4, CipherErrorVecGen_XORInst_1_3_n4,
         CipherErrorVecGen_XORInst_2_3_n4, CipherErrorVecGen_XORInst_3_3_n4,
         CipherErrorVecGen_XORInst_4_3_n4, CipherErrorVecGen_XORInst_5_3_n4,
         CipherErrorVecGen_XORInst_6_3_n4, CipherErrorVecGen_XORInst_7_3_n4,
         CipherErrorVecGen_XORInst_8_3_n4, CipherErrorVecGen_XORInst_9_3_n4,
         CipherErrorVecGen_XORInst_10_3_n4, CipherErrorVecGen_XORInst_11_3_n4,
         CipherErrorVecGen_XORInst_12_3_n4, CipherErrorVecGen_XORInst_13_3_n4,
         CipherErrorVecGen_XORInst_14_3_n4, CipherErrorVecGen_XORInst_15_3_n4,
         SD1_SB_inst_SD1_SB_bit_inst_0_n131,
         SD1_SB_inst_SD1_SB_bit_inst_0_n130,
         SD1_SB_inst_SD1_SB_bit_inst_0_n129,
         SD1_SB_inst_SD1_SB_bit_inst_0_n128,
         SD1_SB_inst_SD1_SB_bit_inst_0_n127,
         SD1_SB_inst_SD1_SB_bit_inst_0_n126,
         SD1_SB_inst_SD1_SB_bit_inst_0_n125,
         SD1_SB_inst_SD1_SB_bit_inst_0_n124,
         SD1_SB_inst_SD1_SB_bit_inst_0_n123,
         SD1_SB_inst_SD1_SB_bit_inst_0_n122,
         SD1_SB_inst_SD1_SB_bit_inst_0_n121,
         SD1_SB_inst_SD1_SB_bit_inst_0_n120,
         SD1_SB_inst_SD1_SB_bit_inst_0_n119,
         SD1_SB_inst_SD1_SB_bit_inst_0_n118,
         SD1_SB_inst_SD1_SB_bit_inst_0_n117,
         SD1_SB_inst_SD1_SB_bit_inst_0_n116,
         SD1_SB_inst_SD1_SB_bit_inst_0_n115,
         SD1_SB_inst_SD1_SB_bit_inst_0_n114,
         SD1_SB_inst_SD1_SB_bit_inst_0_n113,
         SD1_SB_inst_SD1_SB_bit_inst_0_n112,
         SD1_SB_inst_SD1_SB_bit_inst_0_n111,
         SD1_SB_inst_SD1_SB_bit_inst_0_n110,
         SD1_SB_inst_SD1_SB_bit_inst_0_n109,
         SD1_SB_inst_SD1_SB_bit_inst_0_n108,
         SD1_SB_inst_SD1_SB_bit_inst_0_n107,
         SD1_SB_inst_SD1_SB_bit_inst_0_n106,
         SD1_SB_inst_SD1_SB_bit_inst_0_n105,
         SD1_SB_inst_SD1_SB_bit_inst_0_n104,
         SD1_SB_inst_SD1_SB_bit_inst_0_n103,
         SD1_SB_inst_SD1_SB_bit_inst_0_n102,
         SD1_SB_inst_SD1_SB_bit_inst_0_n101,
         SD1_SB_inst_SD1_SB_bit_inst_0_n100, SD1_SB_inst_SD1_SB_bit_inst_0_n99,
         SD1_SB_inst_SD1_SB_bit_inst_0_n98, SD1_SB_inst_SD1_SB_bit_inst_0_n97,
         SD1_SB_inst_SD1_SB_bit_inst_0_n96, SD1_SB_inst_SD1_SB_bit_inst_0_n95,
         SD1_SB_inst_SD1_SB_bit_inst_0_n94, SD1_SB_inst_SD1_SB_bit_inst_0_n93,
         SD1_SB_inst_SD1_SB_bit_inst_0_n92, SD1_SB_inst_SD1_SB_bit_inst_1_n110,
         SD1_SB_inst_SD1_SB_bit_inst_1_n109,
         SD1_SB_inst_SD1_SB_bit_inst_1_n108,
         SD1_SB_inst_SD1_SB_bit_inst_1_n107,
         SD1_SB_inst_SD1_SB_bit_inst_1_n106,
         SD1_SB_inst_SD1_SB_bit_inst_1_n105,
         SD1_SB_inst_SD1_SB_bit_inst_1_n104,
         SD1_SB_inst_SD1_SB_bit_inst_1_n103,
         SD1_SB_inst_SD1_SB_bit_inst_1_n102,
         SD1_SB_inst_SD1_SB_bit_inst_1_n101,
         SD1_SB_inst_SD1_SB_bit_inst_1_n100, SD1_SB_inst_SD1_SB_bit_inst_1_n99,
         SD1_SB_inst_SD1_SB_bit_inst_1_n98, SD1_SB_inst_SD1_SB_bit_inst_1_n97,
         SD1_SB_inst_SD1_SB_bit_inst_1_n96, SD1_SB_inst_SD1_SB_bit_inst_1_n95,
         SD1_SB_inst_SD1_SB_bit_inst_1_n94, SD1_SB_inst_SD1_SB_bit_inst_1_n93,
         SD1_SB_inst_SD1_SB_bit_inst_1_n92, SD1_SB_inst_SD1_SB_bit_inst_1_n91,
         SD1_SB_inst_SD1_SB_bit_inst_1_n90, SD1_SB_inst_SD1_SB_bit_inst_1_n89,
         SD1_SB_inst_SD1_SB_bit_inst_1_n88, SD1_SB_inst_SD1_SB_bit_inst_1_n87,
         SD1_SB_inst_SD1_SB_bit_inst_1_n86, SD1_SB_inst_SD1_SB_bit_inst_1_n85,
         SD1_SB_inst_SD1_SB_bit_inst_1_n84, SD1_SB_inst_SD1_SB_bit_inst_1_n83,
         SD1_SB_inst_SD1_SB_bit_inst_1_n82, SD1_SB_inst_SD1_SB_bit_inst_1_n81,
         SD1_SB_inst_SD1_SB_bit_inst_1_n80, SD1_SB_inst_SD1_SB_bit_inst_1_n79,
         SD1_SB_inst_SD1_SB_bit_inst_1_n78, SD1_SB_inst_SD1_SB_bit_inst_1_n77,
         SD1_SB_inst_SD1_SB_bit_inst_2_n138,
         SD1_SB_inst_SD1_SB_bit_inst_2_n137,
         SD1_SB_inst_SD1_SB_bit_inst_2_n136,
         SD1_SB_inst_SD1_SB_bit_inst_2_n135,
         SD1_SB_inst_SD1_SB_bit_inst_2_n134,
         SD1_SB_inst_SD1_SB_bit_inst_2_n133,
         SD1_SB_inst_SD1_SB_bit_inst_2_n132,
         SD1_SB_inst_SD1_SB_bit_inst_2_n131,
         SD1_SB_inst_SD1_SB_bit_inst_2_n130,
         SD1_SB_inst_SD1_SB_bit_inst_2_n129,
         SD1_SB_inst_SD1_SB_bit_inst_2_n128,
         SD1_SB_inst_SD1_SB_bit_inst_2_n127,
         SD1_SB_inst_SD1_SB_bit_inst_2_n126,
         SD1_SB_inst_SD1_SB_bit_inst_2_n125,
         SD1_SB_inst_SD1_SB_bit_inst_2_n124,
         SD1_SB_inst_SD1_SB_bit_inst_2_n123,
         SD1_SB_inst_SD1_SB_bit_inst_2_n122,
         SD1_SB_inst_SD1_SB_bit_inst_2_n121,
         SD1_SB_inst_SD1_SB_bit_inst_2_n120,
         SD1_SB_inst_SD1_SB_bit_inst_2_n119,
         SD1_SB_inst_SD1_SB_bit_inst_2_n118,
         SD1_SB_inst_SD1_SB_bit_inst_2_n117,
         SD1_SB_inst_SD1_SB_bit_inst_2_n116,
         SD1_SB_inst_SD1_SB_bit_inst_2_n115,
         SD1_SB_inst_SD1_SB_bit_inst_2_n114,
         SD1_SB_inst_SD1_SB_bit_inst_2_n113,
         SD1_SB_inst_SD1_SB_bit_inst_2_n112,
         SD1_SB_inst_SD1_SB_bit_inst_2_n111,
         SD1_SB_inst_SD1_SB_bit_inst_2_n110,
         SD1_SB_inst_SD1_SB_bit_inst_2_n109,
         SD1_SB_inst_SD1_SB_bit_inst_2_n108,
         SD1_SB_inst_SD1_SB_bit_inst_2_n107,
         SD1_SB_inst_SD1_SB_bit_inst_2_n106,
         SD1_SB_inst_SD1_SB_bit_inst_2_n105,
         SD1_SB_inst_SD1_SB_bit_inst_2_n104,
         SD1_SB_inst_SD1_SB_bit_inst_2_n103,
         SD1_SB_inst_SD1_SB_bit_inst_2_n102,
         SD1_SB_inst_SD1_SB_bit_inst_2_n101,
         SD1_SB_inst_SD1_SB_bit_inst_2_n100, SD1_SB_inst_SD1_SB_bit_inst_2_n99,
         SD1_SB_inst_SD1_SB_bit_inst_2_n98, SD1_SB_inst_SD1_SB_bit_inst_2_n97,
         SD1_SB_inst_SD1_SB_bit_inst_3_n141,
         SD1_SB_inst_SD1_SB_bit_inst_3_n140,
         SD1_SB_inst_SD1_SB_bit_inst_3_n139,
         SD1_SB_inst_SD1_SB_bit_inst_3_n138,
         SD1_SB_inst_SD1_SB_bit_inst_3_n137,
         SD1_SB_inst_SD1_SB_bit_inst_3_n136,
         SD1_SB_inst_SD1_SB_bit_inst_3_n135,
         SD1_SB_inst_SD1_SB_bit_inst_3_n134,
         SD1_SB_inst_SD1_SB_bit_inst_3_n133,
         SD1_SB_inst_SD1_SB_bit_inst_3_n132,
         SD1_SB_inst_SD1_SB_bit_inst_3_n131,
         SD1_SB_inst_SD1_SB_bit_inst_3_n130,
         SD1_SB_inst_SD1_SB_bit_inst_3_n129,
         SD1_SB_inst_SD1_SB_bit_inst_3_n128,
         SD1_SB_inst_SD1_SB_bit_inst_3_n127,
         SD1_SB_inst_SD1_SB_bit_inst_3_n126,
         SD1_SB_inst_SD1_SB_bit_inst_3_n125,
         SD1_SB_inst_SD1_SB_bit_inst_3_n124,
         SD1_SB_inst_SD1_SB_bit_inst_3_n123,
         SD1_SB_inst_SD1_SB_bit_inst_3_n122,
         SD1_SB_inst_SD1_SB_bit_inst_3_n121,
         SD1_SB_inst_SD1_SB_bit_inst_3_n120,
         SD1_SB_inst_SD1_SB_bit_inst_3_n119,
         SD1_SB_inst_SD1_SB_bit_inst_3_n118,
         SD1_SB_inst_SD1_SB_bit_inst_3_n117,
         SD1_SB_inst_SD1_SB_bit_inst_3_n116,
         SD1_SB_inst_SD1_SB_bit_inst_3_n115,
         SD1_SB_inst_SD1_SB_bit_inst_3_n114,
         SD1_SB_inst_SD1_SB_bit_inst_3_n113,
         SD1_SB_inst_SD1_SB_bit_inst_3_n112,
         SD1_SB_inst_SD1_SB_bit_inst_3_n111,
         SD1_SB_inst_SD1_SB_bit_inst_3_n110,
         SD1_SB_inst_SD1_SB_bit_inst_3_n109,
         SD1_SB_inst_SD1_SB_bit_inst_3_n108,
         SD1_SB_inst_SD1_SB_bit_inst_3_n107,
         SD1_SB_inst_SD1_SB_bit_inst_3_n106,
         SD1_SB_inst_SD1_SB_bit_inst_3_n105,
         SD1_SB_inst_SD1_SB_bit_inst_3_n104,
         SD1_SB_inst_SD1_SB_bit_inst_3_n103,
         SD1_SB_inst_SD1_SB_bit_inst_3_n102,
         SD1_SB_inst_SD1_SB_bit_inst_3_n101,
         SD1_SB_inst_SD1_SB_bit_inst_3_n100,
         SD1_SB_inst_SD1_SB_bit_inst_4_n131,
         SD1_SB_inst_SD1_SB_bit_inst_4_n130,
         SD1_SB_inst_SD1_SB_bit_inst_4_n129,
         SD1_SB_inst_SD1_SB_bit_inst_4_n128,
         SD1_SB_inst_SD1_SB_bit_inst_4_n127,
         SD1_SB_inst_SD1_SB_bit_inst_4_n126,
         SD1_SB_inst_SD1_SB_bit_inst_4_n125,
         SD1_SB_inst_SD1_SB_bit_inst_4_n124,
         SD1_SB_inst_SD1_SB_bit_inst_4_n123,
         SD1_SB_inst_SD1_SB_bit_inst_4_n122,
         SD1_SB_inst_SD1_SB_bit_inst_4_n121,
         SD1_SB_inst_SD1_SB_bit_inst_4_n120,
         SD1_SB_inst_SD1_SB_bit_inst_4_n119,
         SD1_SB_inst_SD1_SB_bit_inst_4_n118,
         SD1_SB_inst_SD1_SB_bit_inst_4_n117,
         SD1_SB_inst_SD1_SB_bit_inst_4_n116,
         SD1_SB_inst_SD1_SB_bit_inst_4_n115,
         SD1_SB_inst_SD1_SB_bit_inst_4_n114,
         SD1_SB_inst_SD1_SB_bit_inst_4_n113,
         SD1_SB_inst_SD1_SB_bit_inst_4_n112,
         SD1_SB_inst_SD1_SB_bit_inst_4_n111,
         SD1_SB_inst_SD1_SB_bit_inst_4_n110,
         SD1_SB_inst_SD1_SB_bit_inst_4_n109,
         SD1_SB_inst_SD1_SB_bit_inst_4_n108,
         SD1_SB_inst_SD1_SB_bit_inst_4_n107,
         SD1_SB_inst_SD1_SB_bit_inst_4_n106,
         SD1_SB_inst_SD1_SB_bit_inst_4_n105,
         SD1_SB_inst_SD1_SB_bit_inst_4_n104,
         SD1_SB_inst_SD1_SB_bit_inst_4_n103,
         SD1_SB_inst_SD1_SB_bit_inst_4_n102,
         SD1_SB_inst_SD1_SB_bit_inst_4_n101,
         SD1_SB_inst_SD1_SB_bit_inst_4_n100, SD1_SB_inst_SD1_SB_bit_inst_4_n99,
         SD1_SB_inst_SD1_SB_bit_inst_4_n98, SD1_SB_inst_SD1_SB_bit_inst_4_n97,
         SD1_SB_inst_SD1_SB_bit_inst_4_n96, SD1_SB_inst_SD1_SB_bit_inst_4_n95,
         SD1_SB_inst_SD1_SB_bit_inst_4_n94, SD1_SB_inst_SD1_SB_bit_inst_4_n93,
         SD1_SB_inst_SD1_SB_bit_inst_4_n92, SD1_SB_inst_SD1_SB_bit_inst_5_n110,
         SD1_SB_inst_SD1_SB_bit_inst_5_n109,
         SD1_SB_inst_SD1_SB_bit_inst_5_n108,
         SD1_SB_inst_SD1_SB_bit_inst_5_n107,
         SD1_SB_inst_SD1_SB_bit_inst_5_n106,
         SD1_SB_inst_SD1_SB_bit_inst_5_n105,
         SD1_SB_inst_SD1_SB_bit_inst_5_n104,
         SD1_SB_inst_SD1_SB_bit_inst_5_n103,
         SD1_SB_inst_SD1_SB_bit_inst_5_n102,
         SD1_SB_inst_SD1_SB_bit_inst_5_n101,
         SD1_SB_inst_SD1_SB_bit_inst_5_n100, SD1_SB_inst_SD1_SB_bit_inst_5_n99,
         SD1_SB_inst_SD1_SB_bit_inst_5_n98, SD1_SB_inst_SD1_SB_bit_inst_5_n97,
         SD1_SB_inst_SD1_SB_bit_inst_5_n96, SD1_SB_inst_SD1_SB_bit_inst_5_n95,
         SD1_SB_inst_SD1_SB_bit_inst_5_n94, SD1_SB_inst_SD1_SB_bit_inst_5_n93,
         SD1_SB_inst_SD1_SB_bit_inst_5_n92, SD1_SB_inst_SD1_SB_bit_inst_5_n91,
         SD1_SB_inst_SD1_SB_bit_inst_5_n90, SD1_SB_inst_SD1_SB_bit_inst_5_n89,
         SD1_SB_inst_SD1_SB_bit_inst_5_n88, SD1_SB_inst_SD1_SB_bit_inst_5_n87,
         SD1_SB_inst_SD1_SB_bit_inst_5_n86, SD1_SB_inst_SD1_SB_bit_inst_5_n85,
         SD1_SB_inst_SD1_SB_bit_inst_5_n84, SD1_SB_inst_SD1_SB_bit_inst_5_n83,
         SD1_SB_inst_SD1_SB_bit_inst_5_n82, SD1_SB_inst_SD1_SB_bit_inst_5_n81,
         SD1_SB_inst_SD1_SB_bit_inst_5_n80, SD1_SB_inst_SD1_SB_bit_inst_5_n79,
         SD1_SB_inst_SD1_SB_bit_inst_5_n78, SD1_SB_inst_SD1_SB_bit_inst_5_n77,
         SD1_SB_inst_SD1_SB_bit_inst_6_n138,
         SD1_SB_inst_SD1_SB_bit_inst_6_n137,
         SD1_SB_inst_SD1_SB_bit_inst_6_n136,
         SD1_SB_inst_SD1_SB_bit_inst_6_n135,
         SD1_SB_inst_SD1_SB_bit_inst_6_n134,
         SD1_SB_inst_SD1_SB_bit_inst_6_n133,
         SD1_SB_inst_SD1_SB_bit_inst_6_n132,
         SD1_SB_inst_SD1_SB_bit_inst_6_n131,
         SD1_SB_inst_SD1_SB_bit_inst_6_n130,
         SD1_SB_inst_SD1_SB_bit_inst_6_n129,
         SD1_SB_inst_SD1_SB_bit_inst_6_n128,
         SD1_SB_inst_SD1_SB_bit_inst_6_n127,
         SD1_SB_inst_SD1_SB_bit_inst_6_n126,
         SD1_SB_inst_SD1_SB_bit_inst_6_n125,
         SD1_SB_inst_SD1_SB_bit_inst_6_n124,
         SD1_SB_inst_SD1_SB_bit_inst_6_n123,
         SD1_SB_inst_SD1_SB_bit_inst_6_n122,
         SD1_SB_inst_SD1_SB_bit_inst_6_n121,
         SD1_SB_inst_SD1_SB_bit_inst_6_n120,
         SD1_SB_inst_SD1_SB_bit_inst_6_n119,
         SD1_SB_inst_SD1_SB_bit_inst_6_n118,
         SD1_SB_inst_SD1_SB_bit_inst_6_n117,
         SD1_SB_inst_SD1_SB_bit_inst_6_n116,
         SD1_SB_inst_SD1_SB_bit_inst_6_n115,
         SD1_SB_inst_SD1_SB_bit_inst_6_n114,
         SD1_SB_inst_SD1_SB_bit_inst_6_n113,
         SD1_SB_inst_SD1_SB_bit_inst_6_n112,
         SD1_SB_inst_SD1_SB_bit_inst_6_n111,
         SD1_SB_inst_SD1_SB_bit_inst_6_n110,
         SD1_SB_inst_SD1_SB_bit_inst_6_n109,
         SD1_SB_inst_SD1_SB_bit_inst_6_n108,
         SD1_SB_inst_SD1_SB_bit_inst_6_n107,
         SD1_SB_inst_SD1_SB_bit_inst_6_n106,
         SD1_SB_inst_SD1_SB_bit_inst_6_n105,
         SD1_SB_inst_SD1_SB_bit_inst_6_n104,
         SD1_SB_inst_SD1_SB_bit_inst_6_n103,
         SD1_SB_inst_SD1_SB_bit_inst_6_n102,
         SD1_SB_inst_SD1_SB_bit_inst_6_n101,
         SD1_SB_inst_SD1_SB_bit_inst_6_n100, SD1_SB_inst_SD1_SB_bit_inst_6_n99,
         SD1_SB_inst_SD1_SB_bit_inst_6_n98, SD1_SB_inst_SD1_SB_bit_inst_6_n97,
         SD1_SB_inst_SD1_SB_bit_inst_7_n141,
         SD1_SB_inst_SD1_SB_bit_inst_7_n140,
         SD1_SB_inst_SD1_SB_bit_inst_7_n139,
         SD1_SB_inst_SD1_SB_bit_inst_7_n138,
         SD1_SB_inst_SD1_SB_bit_inst_7_n137,
         SD1_SB_inst_SD1_SB_bit_inst_7_n136,
         SD1_SB_inst_SD1_SB_bit_inst_7_n135,
         SD1_SB_inst_SD1_SB_bit_inst_7_n134,
         SD1_SB_inst_SD1_SB_bit_inst_7_n133,
         SD1_SB_inst_SD1_SB_bit_inst_7_n132,
         SD1_SB_inst_SD1_SB_bit_inst_7_n131,
         SD1_SB_inst_SD1_SB_bit_inst_7_n130,
         SD1_SB_inst_SD1_SB_bit_inst_7_n129,
         SD1_SB_inst_SD1_SB_bit_inst_7_n128,
         SD1_SB_inst_SD1_SB_bit_inst_7_n127,
         SD1_SB_inst_SD1_SB_bit_inst_7_n126,
         SD1_SB_inst_SD1_SB_bit_inst_7_n125,
         SD1_SB_inst_SD1_SB_bit_inst_7_n124,
         SD1_SB_inst_SD1_SB_bit_inst_7_n123,
         SD1_SB_inst_SD1_SB_bit_inst_7_n122,
         SD1_SB_inst_SD1_SB_bit_inst_7_n121,
         SD1_SB_inst_SD1_SB_bit_inst_7_n120,
         SD1_SB_inst_SD1_SB_bit_inst_7_n119,
         SD1_SB_inst_SD1_SB_bit_inst_7_n118,
         SD1_SB_inst_SD1_SB_bit_inst_7_n117,
         SD1_SB_inst_SD1_SB_bit_inst_7_n116,
         SD1_SB_inst_SD1_SB_bit_inst_7_n115,
         SD1_SB_inst_SD1_SB_bit_inst_7_n114,
         SD1_SB_inst_SD1_SB_bit_inst_7_n113,
         SD1_SB_inst_SD1_SB_bit_inst_7_n112,
         SD1_SB_inst_SD1_SB_bit_inst_7_n111,
         SD1_SB_inst_SD1_SB_bit_inst_7_n110,
         SD1_SB_inst_SD1_SB_bit_inst_7_n109,
         SD1_SB_inst_SD1_SB_bit_inst_7_n108,
         SD1_SB_inst_SD1_SB_bit_inst_7_n107,
         SD1_SB_inst_SD1_SB_bit_inst_7_n106,
         SD1_SB_inst_SD1_SB_bit_inst_7_n105,
         SD1_SB_inst_SD1_SB_bit_inst_7_n104,
         SD1_SB_inst_SD1_SB_bit_inst_7_n103,
         SD1_SB_inst_SD1_SB_bit_inst_7_n102,
         SD1_SB_inst_SD1_SB_bit_inst_7_n101,
         SD1_SB_inst_SD1_SB_bit_inst_7_n100,
         SD1_SB_inst_SD1_SB_bit_inst_8_n131,
         SD1_SB_inst_SD1_SB_bit_inst_8_n130,
         SD1_SB_inst_SD1_SB_bit_inst_8_n129,
         SD1_SB_inst_SD1_SB_bit_inst_8_n128,
         SD1_SB_inst_SD1_SB_bit_inst_8_n127,
         SD1_SB_inst_SD1_SB_bit_inst_8_n126,
         SD1_SB_inst_SD1_SB_bit_inst_8_n125,
         SD1_SB_inst_SD1_SB_bit_inst_8_n124,
         SD1_SB_inst_SD1_SB_bit_inst_8_n123,
         SD1_SB_inst_SD1_SB_bit_inst_8_n122,
         SD1_SB_inst_SD1_SB_bit_inst_8_n121,
         SD1_SB_inst_SD1_SB_bit_inst_8_n120,
         SD1_SB_inst_SD1_SB_bit_inst_8_n119,
         SD1_SB_inst_SD1_SB_bit_inst_8_n118,
         SD1_SB_inst_SD1_SB_bit_inst_8_n117,
         SD1_SB_inst_SD1_SB_bit_inst_8_n116,
         SD1_SB_inst_SD1_SB_bit_inst_8_n115,
         SD1_SB_inst_SD1_SB_bit_inst_8_n114,
         SD1_SB_inst_SD1_SB_bit_inst_8_n113,
         SD1_SB_inst_SD1_SB_bit_inst_8_n112,
         SD1_SB_inst_SD1_SB_bit_inst_8_n111,
         SD1_SB_inst_SD1_SB_bit_inst_8_n110,
         SD1_SB_inst_SD1_SB_bit_inst_8_n109,
         SD1_SB_inst_SD1_SB_bit_inst_8_n108,
         SD1_SB_inst_SD1_SB_bit_inst_8_n107,
         SD1_SB_inst_SD1_SB_bit_inst_8_n106,
         SD1_SB_inst_SD1_SB_bit_inst_8_n105,
         SD1_SB_inst_SD1_SB_bit_inst_8_n104,
         SD1_SB_inst_SD1_SB_bit_inst_8_n103,
         SD1_SB_inst_SD1_SB_bit_inst_8_n102,
         SD1_SB_inst_SD1_SB_bit_inst_8_n101,
         SD1_SB_inst_SD1_SB_bit_inst_8_n100, SD1_SB_inst_SD1_SB_bit_inst_8_n99,
         SD1_SB_inst_SD1_SB_bit_inst_8_n98, SD1_SB_inst_SD1_SB_bit_inst_8_n97,
         SD1_SB_inst_SD1_SB_bit_inst_8_n96, SD1_SB_inst_SD1_SB_bit_inst_8_n95,
         SD1_SB_inst_SD1_SB_bit_inst_8_n94, SD1_SB_inst_SD1_SB_bit_inst_8_n93,
         SD1_SB_inst_SD1_SB_bit_inst_8_n92, SD1_SB_inst_SD1_SB_bit_inst_9_n110,
         SD1_SB_inst_SD1_SB_bit_inst_9_n109,
         SD1_SB_inst_SD1_SB_bit_inst_9_n108,
         SD1_SB_inst_SD1_SB_bit_inst_9_n107,
         SD1_SB_inst_SD1_SB_bit_inst_9_n106,
         SD1_SB_inst_SD1_SB_bit_inst_9_n105,
         SD1_SB_inst_SD1_SB_bit_inst_9_n104,
         SD1_SB_inst_SD1_SB_bit_inst_9_n103,
         SD1_SB_inst_SD1_SB_bit_inst_9_n102,
         SD1_SB_inst_SD1_SB_bit_inst_9_n101,
         SD1_SB_inst_SD1_SB_bit_inst_9_n100, SD1_SB_inst_SD1_SB_bit_inst_9_n99,
         SD1_SB_inst_SD1_SB_bit_inst_9_n98, SD1_SB_inst_SD1_SB_bit_inst_9_n97,
         SD1_SB_inst_SD1_SB_bit_inst_9_n96, SD1_SB_inst_SD1_SB_bit_inst_9_n95,
         SD1_SB_inst_SD1_SB_bit_inst_9_n94, SD1_SB_inst_SD1_SB_bit_inst_9_n93,
         SD1_SB_inst_SD1_SB_bit_inst_9_n92, SD1_SB_inst_SD1_SB_bit_inst_9_n91,
         SD1_SB_inst_SD1_SB_bit_inst_9_n90, SD1_SB_inst_SD1_SB_bit_inst_9_n89,
         SD1_SB_inst_SD1_SB_bit_inst_9_n88, SD1_SB_inst_SD1_SB_bit_inst_9_n87,
         SD1_SB_inst_SD1_SB_bit_inst_9_n86, SD1_SB_inst_SD1_SB_bit_inst_9_n85,
         SD1_SB_inst_SD1_SB_bit_inst_9_n84, SD1_SB_inst_SD1_SB_bit_inst_9_n83,
         SD1_SB_inst_SD1_SB_bit_inst_9_n82, SD1_SB_inst_SD1_SB_bit_inst_9_n81,
         SD1_SB_inst_SD1_SB_bit_inst_9_n80, SD1_SB_inst_SD1_SB_bit_inst_9_n79,
         SD1_SB_inst_SD1_SB_bit_inst_9_n78, SD1_SB_inst_SD1_SB_bit_inst_9_n77,
         SD1_SB_inst_SD1_SB_bit_inst_10_n138,
         SD1_SB_inst_SD1_SB_bit_inst_10_n137,
         SD1_SB_inst_SD1_SB_bit_inst_10_n136,
         SD1_SB_inst_SD1_SB_bit_inst_10_n135,
         SD1_SB_inst_SD1_SB_bit_inst_10_n134,
         SD1_SB_inst_SD1_SB_bit_inst_10_n133,
         SD1_SB_inst_SD1_SB_bit_inst_10_n132,
         SD1_SB_inst_SD1_SB_bit_inst_10_n131,
         SD1_SB_inst_SD1_SB_bit_inst_10_n130,
         SD1_SB_inst_SD1_SB_bit_inst_10_n129,
         SD1_SB_inst_SD1_SB_bit_inst_10_n128,
         SD1_SB_inst_SD1_SB_bit_inst_10_n127,
         SD1_SB_inst_SD1_SB_bit_inst_10_n126,
         SD1_SB_inst_SD1_SB_bit_inst_10_n125,
         SD1_SB_inst_SD1_SB_bit_inst_10_n124,
         SD1_SB_inst_SD1_SB_bit_inst_10_n123,
         SD1_SB_inst_SD1_SB_bit_inst_10_n122,
         SD1_SB_inst_SD1_SB_bit_inst_10_n121,
         SD1_SB_inst_SD1_SB_bit_inst_10_n120,
         SD1_SB_inst_SD1_SB_bit_inst_10_n119,
         SD1_SB_inst_SD1_SB_bit_inst_10_n118,
         SD1_SB_inst_SD1_SB_bit_inst_10_n117,
         SD1_SB_inst_SD1_SB_bit_inst_10_n116,
         SD1_SB_inst_SD1_SB_bit_inst_10_n115,
         SD1_SB_inst_SD1_SB_bit_inst_10_n114,
         SD1_SB_inst_SD1_SB_bit_inst_10_n113,
         SD1_SB_inst_SD1_SB_bit_inst_10_n112,
         SD1_SB_inst_SD1_SB_bit_inst_10_n111,
         SD1_SB_inst_SD1_SB_bit_inst_10_n110,
         SD1_SB_inst_SD1_SB_bit_inst_10_n109,
         SD1_SB_inst_SD1_SB_bit_inst_10_n108,
         SD1_SB_inst_SD1_SB_bit_inst_10_n107,
         SD1_SB_inst_SD1_SB_bit_inst_10_n106,
         SD1_SB_inst_SD1_SB_bit_inst_10_n105,
         SD1_SB_inst_SD1_SB_bit_inst_10_n104,
         SD1_SB_inst_SD1_SB_bit_inst_10_n103,
         SD1_SB_inst_SD1_SB_bit_inst_10_n102,
         SD1_SB_inst_SD1_SB_bit_inst_10_n101,
         SD1_SB_inst_SD1_SB_bit_inst_10_n100,
         SD1_SB_inst_SD1_SB_bit_inst_10_n99,
         SD1_SB_inst_SD1_SB_bit_inst_10_n98,
         SD1_SB_inst_SD1_SB_bit_inst_10_n97,
         SD1_SB_inst_SD1_SB_bit_inst_11_n141,
         SD1_SB_inst_SD1_SB_bit_inst_11_n140,
         SD1_SB_inst_SD1_SB_bit_inst_11_n139,
         SD1_SB_inst_SD1_SB_bit_inst_11_n138,
         SD1_SB_inst_SD1_SB_bit_inst_11_n137,
         SD1_SB_inst_SD1_SB_bit_inst_11_n136,
         SD1_SB_inst_SD1_SB_bit_inst_11_n135,
         SD1_SB_inst_SD1_SB_bit_inst_11_n134,
         SD1_SB_inst_SD1_SB_bit_inst_11_n133,
         SD1_SB_inst_SD1_SB_bit_inst_11_n132,
         SD1_SB_inst_SD1_SB_bit_inst_11_n131,
         SD1_SB_inst_SD1_SB_bit_inst_11_n130,
         SD1_SB_inst_SD1_SB_bit_inst_11_n129,
         SD1_SB_inst_SD1_SB_bit_inst_11_n128,
         SD1_SB_inst_SD1_SB_bit_inst_11_n127,
         SD1_SB_inst_SD1_SB_bit_inst_11_n126,
         SD1_SB_inst_SD1_SB_bit_inst_11_n125,
         SD1_SB_inst_SD1_SB_bit_inst_11_n124,
         SD1_SB_inst_SD1_SB_bit_inst_11_n123,
         SD1_SB_inst_SD1_SB_bit_inst_11_n122,
         SD1_SB_inst_SD1_SB_bit_inst_11_n121,
         SD1_SB_inst_SD1_SB_bit_inst_11_n120,
         SD1_SB_inst_SD1_SB_bit_inst_11_n119,
         SD1_SB_inst_SD1_SB_bit_inst_11_n118,
         SD1_SB_inst_SD1_SB_bit_inst_11_n117,
         SD1_SB_inst_SD1_SB_bit_inst_11_n116,
         SD1_SB_inst_SD1_SB_bit_inst_11_n115,
         SD1_SB_inst_SD1_SB_bit_inst_11_n114,
         SD1_SB_inst_SD1_SB_bit_inst_11_n113,
         SD1_SB_inst_SD1_SB_bit_inst_11_n112,
         SD1_SB_inst_SD1_SB_bit_inst_11_n111,
         SD1_SB_inst_SD1_SB_bit_inst_11_n110,
         SD1_SB_inst_SD1_SB_bit_inst_11_n109,
         SD1_SB_inst_SD1_SB_bit_inst_11_n108,
         SD1_SB_inst_SD1_SB_bit_inst_11_n107,
         SD1_SB_inst_SD1_SB_bit_inst_11_n106,
         SD1_SB_inst_SD1_SB_bit_inst_11_n105,
         SD1_SB_inst_SD1_SB_bit_inst_11_n104,
         SD1_SB_inst_SD1_SB_bit_inst_11_n103,
         SD1_SB_inst_SD1_SB_bit_inst_11_n102,
         SD1_SB_inst_SD1_SB_bit_inst_11_n101,
         SD1_SB_inst_SD1_SB_bit_inst_11_n100,
         SD1_SB_inst_SD1_SB_bit_inst_12_n131,
         SD1_SB_inst_SD1_SB_bit_inst_12_n130,
         SD1_SB_inst_SD1_SB_bit_inst_12_n129,
         SD1_SB_inst_SD1_SB_bit_inst_12_n128,
         SD1_SB_inst_SD1_SB_bit_inst_12_n127,
         SD1_SB_inst_SD1_SB_bit_inst_12_n126,
         SD1_SB_inst_SD1_SB_bit_inst_12_n125,
         SD1_SB_inst_SD1_SB_bit_inst_12_n124,
         SD1_SB_inst_SD1_SB_bit_inst_12_n123,
         SD1_SB_inst_SD1_SB_bit_inst_12_n122,
         SD1_SB_inst_SD1_SB_bit_inst_12_n121,
         SD1_SB_inst_SD1_SB_bit_inst_12_n120,
         SD1_SB_inst_SD1_SB_bit_inst_12_n119,
         SD1_SB_inst_SD1_SB_bit_inst_12_n118,
         SD1_SB_inst_SD1_SB_bit_inst_12_n117,
         SD1_SB_inst_SD1_SB_bit_inst_12_n116,
         SD1_SB_inst_SD1_SB_bit_inst_12_n115,
         SD1_SB_inst_SD1_SB_bit_inst_12_n114,
         SD1_SB_inst_SD1_SB_bit_inst_12_n113,
         SD1_SB_inst_SD1_SB_bit_inst_12_n112,
         SD1_SB_inst_SD1_SB_bit_inst_12_n111,
         SD1_SB_inst_SD1_SB_bit_inst_12_n110,
         SD1_SB_inst_SD1_SB_bit_inst_12_n109,
         SD1_SB_inst_SD1_SB_bit_inst_12_n108,
         SD1_SB_inst_SD1_SB_bit_inst_12_n107,
         SD1_SB_inst_SD1_SB_bit_inst_12_n106,
         SD1_SB_inst_SD1_SB_bit_inst_12_n105,
         SD1_SB_inst_SD1_SB_bit_inst_12_n104,
         SD1_SB_inst_SD1_SB_bit_inst_12_n103,
         SD1_SB_inst_SD1_SB_bit_inst_12_n102,
         SD1_SB_inst_SD1_SB_bit_inst_12_n101,
         SD1_SB_inst_SD1_SB_bit_inst_12_n100,
         SD1_SB_inst_SD1_SB_bit_inst_12_n99,
         SD1_SB_inst_SD1_SB_bit_inst_12_n98,
         SD1_SB_inst_SD1_SB_bit_inst_12_n97,
         SD1_SB_inst_SD1_SB_bit_inst_12_n96,
         SD1_SB_inst_SD1_SB_bit_inst_12_n95,
         SD1_SB_inst_SD1_SB_bit_inst_12_n94,
         SD1_SB_inst_SD1_SB_bit_inst_12_n93,
         SD1_SB_inst_SD1_SB_bit_inst_12_n92,
         SD1_SB_inst_SD1_SB_bit_inst_13_n110,
         SD1_SB_inst_SD1_SB_bit_inst_13_n109,
         SD1_SB_inst_SD1_SB_bit_inst_13_n108,
         SD1_SB_inst_SD1_SB_bit_inst_13_n107,
         SD1_SB_inst_SD1_SB_bit_inst_13_n106,
         SD1_SB_inst_SD1_SB_bit_inst_13_n105,
         SD1_SB_inst_SD1_SB_bit_inst_13_n104,
         SD1_SB_inst_SD1_SB_bit_inst_13_n103,
         SD1_SB_inst_SD1_SB_bit_inst_13_n102,
         SD1_SB_inst_SD1_SB_bit_inst_13_n101,
         SD1_SB_inst_SD1_SB_bit_inst_13_n100,
         SD1_SB_inst_SD1_SB_bit_inst_13_n99,
         SD1_SB_inst_SD1_SB_bit_inst_13_n98,
         SD1_SB_inst_SD1_SB_bit_inst_13_n97,
         SD1_SB_inst_SD1_SB_bit_inst_13_n96,
         SD1_SB_inst_SD1_SB_bit_inst_13_n95,
         SD1_SB_inst_SD1_SB_bit_inst_13_n94,
         SD1_SB_inst_SD1_SB_bit_inst_13_n93,
         SD1_SB_inst_SD1_SB_bit_inst_13_n92,
         SD1_SB_inst_SD1_SB_bit_inst_13_n91,
         SD1_SB_inst_SD1_SB_bit_inst_13_n90,
         SD1_SB_inst_SD1_SB_bit_inst_13_n89,
         SD1_SB_inst_SD1_SB_bit_inst_13_n88,
         SD1_SB_inst_SD1_SB_bit_inst_13_n87,
         SD1_SB_inst_SD1_SB_bit_inst_13_n86,
         SD1_SB_inst_SD1_SB_bit_inst_13_n85,
         SD1_SB_inst_SD1_SB_bit_inst_13_n84,
         SD1_SB_inst_SD1_SB_bit_inst_13_n83,
         SD1_SB_inst_SD1_SB_bit_inst_13_n82,
         SD1_SB_inst_SD1_SB_bit_inst_13_n81,
         SD1_SB_inst_SD1_SB_bit_inst_13_n80,
         SD1_SB_inst_SD1_SB_bit_inst_13_n79,
         SD1_SB_inst_SD1_SB_bit_inst_13_n78,
         SD1_SB_inst_SD1_SB_bit_inst_13_n77,
         SD1_SB_inst_SD1_SB_bit_inst_14_n138,
         SD1_SB_inst_SD1_SB_bit_inst_14_n137,
         SD1_SB_inst_SD1_SB_bit_inst_14_n136,
         SD1_SB_inst_SD1_SB_bit_inst_14_n135,
         SD1_SB_inst_SD1_SB_bit_inst_14_n134,
         SD1_SB_inst_SD1_SB_bit_inst_14_n133,
         SD1_SB_inst_SD1_SB_bit_inst_14_n132,
         SD1_SB_inst_SD1_SB_bit_inst_14_n131,
         SD1_SB_inst_SD1_SB_bit_inst_14_n130,
         SD1_SB_inst_SD1_SB_bit_inst_14_n129,
         SD1_SB_inst_SD1_SB_bit_inst_14_n128,
         SD1_SB_inst_SD1_SB_bit_inst_14_n127,
         SD1_SB_inst_SD1_SB_bit_inst_14_n126,
         SD1_SB_inst_SD1_SB_bit_inst_14_n125,
         SD1_SB_inst_SD1_SB_bit_inst_14_n124,
         SD1_SB_inst_SD1_SB_bit_inst_14_n123,
         SD1_SB_inst_SD1_SB_bit_inst_14_n122,
         SD1_SB_inst_SD1_SB_bit_inst_14_n121,
         SD1_SB_inst_SD1_SB_bit_inst_14_n120,
         SD1_SB_inst_SD1_SB_bit_inst_14_n119,
         SD1_SB_inst_SD1_SB_bit_inst_14_n118,
         SD1_SB_inst_SD1_SB_bit_inst_14_n117,
         SD1_SB_inst_SD1_SB_bit_inst_14_n116,
         SD1_SB_inst_SD1_SB_bit_inst_14_n115,
         SD1_SB_inst_SD1_SB_bit_inst_14_n114,
         SD1_SB_inst_SD1_SB_bit_inst_14_n113,
         SD1_SB_inst_SD1_SB_bit_inst_14_n112,
         SD1_SB_inst_SD1_SB_bit_inst_14_n111,
         SD1_SB_inst_SD1_SB_bit_inst_14_n110,
         SD1_SB_inst_SD1_SB_bit_inst_14_n109,
         SD1_SB_inst_SD1_SB_bit_inst_14_n108,
         SD1_SB_inst_SD1_SB_bit_inst_14_n107,
         SD1_SB_inst_SD1_SB_bit_inst_14_n106,
         SD1_SB_inst_SD1_SB_bit_inst_14_n105,
         SD1_SB_inst_SD1_SB_bit_inst_14_n104,
         SD1_SB_inst_SD1_SB_bit_inst_14_n103,
         SD1_SB_inst_SD1_SB_bit_inst_14_n102,
         SD1_SB_inst_SD1_SB_bit_inst_14_n101,
         SD1_SB_inst_SD1_SB_bit_inst_14_n100,
         SD1_SB_inst_SD1_SB_bit_inst_14_n99,
         SD1_SB_inst_SD1_SB_bit_inst_14_n98,
         SD1_SB_inst_SD1_SB_bit_inst_14_n97,
         SD1_SB_inst_SD1_SB_bit_inst_15_n141,
         SD1_SB_inst_SD1_SB_bit_inst_15_n140,
         SD1_SB_inst_SD1_SB_bit_inst_15_n139,
         SD1_SB_inst_SD1_SB_bit_inst_15_n138,
         SD1_SB_inst_SD1_SB_bit_inst_15_n137,
         SD1_SB_inst_SD1_SB_bit_inst_15_n136,
         SD1_SB_inst_SD1_SB_bit_inst_15_n135,
         SD1_SB_inst_SD1_SB_bit_inst_15_n134,
         SD1_SB_inst_SD1_SB_bit_inst_15_n133,
         SD1_SB_inst_SD1_SB_bit_inst_15_n132,
         SD1_SB_inst_SD1_SB_bit_inst_15_n131,
         SD1_SB_inst_SD1_SB_bit_inst_15_n130,
         SD1_SB_inst_SD1_SB_bit_inst_15_n129,
         SD1_SB_inst_SD1_SB_bit_inst_15_n128,
         SD1_SB_inst_SD1_SB_bit_inst_15_n127,
         SD1_SB_inst_SD1_SB_bit_inst_15_n126,
         SD1_SB_inst_SD1_SB_bit_inst_15_n125,
         SD1_SB_inst_SD1_SB_bit_inst_15_n124,
         SD1_SB_inst_SD1_SB_bit_inst_15_n123,
         SD1_SB_inst_SD1_SB_bit_inst_15_n122,
         SD1_SB_inst_SD1_SB_bit_inst_15_n121,
         SD1_SB_inst_SD1_SB_bit_inst_15_n120,
         SD1_SB_inst_SD1_SB_bit_inst_15_n119,
         SD1_SB_inst_SD1_SB_bit_inst_15_n118,
         SD1_SB_inst_SD1_SB_bit_inst_15_n117,
         SD1_SB_inst_SD1_SB_bit_inst_15_n116,
         SD1_SB_inst_SD1_SB_bit_inst_15_n115,
         SD1_SB_inst_SD1_SB_bit_inst_15_n114,
         SD1_SB_inst_SD1_SB_bit_inst_15_n113,
         SD1_SB_inst_SD1_SB_bit_inst_15_n112,
         SD1_SB_inst_SD1_SB_bit_inst_15_n111,
         SD1_SB_inst_SD1_SB_bit_inst_15_n110,
         SD1_SB_inst_SD1_SB_bit_inst_15_n109,
         SD1_SB_inst_SD1_SB_bit_inst_15_n108,
         SD1_SB_inst_SD1_SB_bit_inst_15_n107,
         SD1_SB_inst_SD1_SB_bit_inst_15_n106,
         SD1_SB_inst_SD1_SB_bit_inst_15_n105,
         SD1_SB_inst_SD1_SB_bit_inst_15_n104,
         SD1_SB_inst_SD1_SB_bit_inst_15_n103,
         SD1_SB_inst_SD1_SB_bit_inst_15_n102,
         SD1_SB_inst_SD1_SB_bit_inst_15_n101,
         SD1_SB_inst_SD1_SB_bit_inst_15_n100,
         SD1_SB_inst_SD1_SB_bit_inst_16_n132,
         SD1_SB_inst_SD1_SB_bit_inst_16_n131,
         SD1_SB_inst_SD1_SB_bit_inst_16_n130,
         SD1_SB_inst_SD1_SB_bit_inst_16_n129,
         SD1_SB_inst_SD1_SB_bit_inst_16_n128,
         SD1_SB_inst_SD1_SB_bit_inst_16_n127,
         SD1_SB_inst_SD1_SB_bit_inst_16_n126,
         SD1_SB_inst_SD1_SB_bit_inst_16_n125,
         SD1_SB_inst_SD1_SB_bit_inst_16_n124,
         SD1_SB_inst_SD1_SB_bit_inst_16_n123,
         SD1_SB_inst_SD1_SB_bit_inst_16_n122,
         SD1_SB_inst_SD1_SB_bit_inst_16_n121,
         SD1_SB_inst_SD1_SB_bit_inst_16_n120,
         SD1_SB_inst_SD1_SB_bit_inst_16_n119,
         SD1_SB_inst_SD1_SB_bit_inst_16_n118,
         SD1_SB_inst_SD1_SB_bit_inst_16_n117,
         SD1_SB_inst_SD1_SB_bit_inst_16_n116,
         SD1_SB_inst_SD1_SB_bit_inst_16_n115,
         SD1_SB_inst_SD1_SB_bit_inst_16_n114,
         SD1_SB_inst_SD1_SB_bit_inst_16_n113,
         SD1_SB_inst_SD1_SB_bit_inst_16_n112,
         SD1_SB_inst_SD1_SB_bit_inst_16_n111,
         SD1_SB_inst_SD1_SB_bit_inst_16_n110,
         SD1_SB_inst_SD1_SB_bit_inst_16_n109,
         SD1_SB_inst_SD1_SB_bit_inst_16_n108,
         SD1_SB_inst_SD1_SB_bit_inst_16_n107,
         SD1_SB_inst_SD1_SB_bit_inst_16_n106,
         SD1_SB_inst_SD1_SB_bit_inst_16_n105,
         SD1_SB_inst_SD1_SB_bit_inst_16_n104,
         SD1_SB_inst_SD1_SB_bit_inst_16_n103,
         SD1_SB_inst_SD1_SB_bit_inst_16_n102,
         SD1_SB_inst_SD1_SB_bit_inst_16_n101,
         SD1_SB_inst_SD1_SB_bit_inst_16_n100,
         SD1_SB_inst_SD1_SB_bit_inst_16_n99,
         SD1_SB_inst_SD1_SB_bit_inst_16_n98,
         SD1_SB_inst_SD1_SB_bit_inst_16_n97,
         SD1_SB_inst_SD1_SB_bit_inst_16_n96,
         SD1_SB_inst_SD1_SB_bit_inst_16_n95,
         SD1_SB_inst_SD1_SB_bit_inst_16_n94,
         SD1_SB_inst_SD1_SB_bit_inst_16_n93,
         SD1_SB_inst_SD1_SB_bit_inst_16_n92,
         SD1_SB_inst_SD1_SB_bit_inst_17_n109,
         SD1_SB_inst_SD1_SB_bit_inst_17_n108,
         SD1_SB_inst_SD1_SB_bit_inst_17_n107,
         SD1_SB_inst_SD1_SB_bit_inst_17_n106,
         SD1_SB_inst_SD1_SB_bit_inst_17_n105,
         SD1_SB_inst_SD1_SB_bit_inst_17_n104,
         SD1_SB_inst_SD1_SB_bit_inst_17_n103,
         SD1_SB_inst_SD1_SB_bit_inst_17_n102,
         SD1_SB_inst_SD1_SB_bit_inst_17_n101,
         SD1_SB_inst_SD1_SB_bit_inst_17_n100,
         SD1_SB_inst_SD1_SB_bit_inst_17_n99,
         SD1_SB_inst_SD1_SB_bit_inst_17_n98,
         SD1_SB_inst_SD1_SB_bit_inst_17_n97,
         SD1_SB_inst_SD1_SB_bit_inst_17_n96,
         SD1_SB_inst_SD1_SB_bit_inst_17_n95,
         SD1_SB_inst_SD1_SB_bit_inst_17_n94,
         SD1_SB_inst_SD1_SB_bit_inst_17_n93,
         SD1_SB_inst_SD1_SB_bit_inst_17_n92,
         SD1_SB_inst_SD1_SB_bit_inst_17_n91,
         SD1_SB_inst_SD1_SB_bit_inst_17_n90,
         SD1_SB_inst_SD1_SB_bit_inst_17_n89,
         SD1_SB_inst_SD1_SB_bit_inst_17_n88,
         SD1_SB_inst_SD1_SB_bit_inst_17_n87,
         SD1_SB_inst_SD1_SB_bit_inst_17_n86,
         SD1_SB_inst_SD1_SB_bit_inst_17_n85,
         SD1_SB_inst_SD1_SB_bit_inst_17_n84,
         SD1_SB_inst_SD1_SB_bit_inst_17_n83,
         SD1_SB_inst_SD1_SB_bit_inst_17_n82,
         SD1_SB_inst_SD1_SB_bit_inst_17_n81,
         SD1_SB_inst_SD1_SB_bit_inst_17_n80,
         SD1_SB_inst_SD1_SB_bit_inst_17_n79,
         SD1_SB_inst_SD1_SB_bit_inst_17_n78,
         SD1_SB_inst_SD1_SB_bit_inst_17_n77,
         SD1_SB_inst_SD1_SB_bit_inst_18_n137,
         SD1_SB_inst_SD1_SB_bit_inst_18_n136,
         SD1_SB_inst_SD1_SB_bit_inst_18_n135,
         SD1_SB_inst_SD1_SB_bit_inst_18_n134,
         SD1_SB_inst_SD1_SB_bit_inst_18_n133,
         SD1_SB_inst_SD1_SB_bit_inst_18_n132,
         SD1_SB_inst_SD1_SB_bit_inst_18_n131,
         SD1_SB_inst_SD1_SB_bit_inst_18_n130,
         SD1_SB_inst_SD1_SB_bit_inst_18_n129,
         SD1_SB_inst_SD1_SB_bit_inst_18_n128,
         SD1_SB_inst_SD1_SB_bit_inst_18_n127,
         SD1_SB_inst_SD1_SB_bit_inst_18_n126,
         SD1_SB_inst_SD1_SB_bit_inst_18_n125,
         SD1_SB_inst_SD1_SB_bit_inst_18_n124,
         SD1_SB_inst_SD1_SB_bit_inst_18_n123,
         SD1_SB_inst_SD1_SB_bit_inst_18_n122,
         SD1_SB_inst_SD1_SB_bit_inst_18_n121,
         SD1_SB_inst_SD1_SB_bit_inst_18_n120,
         SD1_SB_inst_SD1_SB_bit_inst_18_n119,
         SD1_SB_inst_SD1_SB_bit_inst_18_n118,
         SD1_SB_inst_SD1_SB_bit_inst_18_n117,
         SD1_SB_inst_SD1_SB_bit_inst_18_n116,
         SD1_SB_inst_SD1_SB_bit_inst_18_n115,
         SD1_SB_inst_SD1_SB_bit_inst_18_n114,
         SD1_SB_inst_SD1_SB_bit_inst_18_n113,
         SD1_SB_inst_SD1_SB_bit_inst_18_n112,
         SD1_SB_inst_SD1_SB_bit_inst_18_n111,
         SD1_SB_inst_SD1_SB_bit_inst_18_n110,
         SD1_SB_inst_SD1_SB_bit_inst_18_n109,
         SD1_SB_inst_SD1_SB_bit_inst_18_n108,
         SD1_SB_inst_SD1_SB_bit_inst_18_n107,
         SD1_SB_inst_SD1_SB_bit_inst_18_n106,
         SD1_SB_inst_SD1_SB_bit_inst_18_n105,
         SD1_SB_inst_SD1_SB_bit_inst_18_n104,
         SD1_SB_inst_SD1_SB_bit_inst_18_n103,
         SD1_SB_inst_SD1_SB_bit_inst_18_n102,
         SD1_SB_inst_SD1_SB_bit_inst_18_n101,
         SD1_SB_inst_SD1_SB_bit_inst_18_n100,
         SD1_SB_inst_SD1_SB_bit_inst_18_n99,
         SD1_SB_inst_SD1_SB_bit_inst_18_n98,
         SD1_SB_inst_SD1_SB_bit_inst_18_n97,
         SD1_SB_inst_SD1_SB_bit_inst_19_n141,
         SD1_SB_inst_SD1_SB_bit_inst_19_n140,
         SD1_SB_inst_SD1_SB_bit_inst_19_n139,
         SD1_SB_inst_SD1_SB_bit_inst_19_n138,
         SD1_SB_inst_SD1_SB_bit_inst_19_n137,
         SD1_SB_inst_SD1_SB_bit_inst_19_n136,
         SD1_SB_inst_SD1_SB_bit_inst_19_n135,
         SD1_SB_inst_SD1_SB_bit_inst_19_n134,
         SD1_SB_inst_SD1_SB_bit_inst_19_n133,
         SD1_SB_inst_SD1_SB_bit_inst_19_n132,
         SD1_SB_inst_SD1_SB_bit_inst_19_n131,
         SD1_SB_inst_SD1_SB_bit_inst_19_n130,
         SD1_SB_inst_SD1_SB_bit_inst_19_n129,
         SD1_SB_inst_SD1_SB_bit_inst_19_n128,
         SD1_SB_inst_SD1_SB_bit_inst_19_n127,
         SD1_SB_inst_SD1_SB_bit_inst_19_n126,
         SD1_SB_inst_SD1_SB_bit_inst_19_n125,
         SD1_SB_inst_SD1_SB_bit_inst_19_n124,
         SD1_SB_inst_SD1_SB_bit_inst_19_n123,
         SD1_SB_inst_SD1_SB_bit_inst_19_n122,
         SD1_SB_inst_SD1_SB_bit_inst_19_n121,
         SD1_SB_inst_SD1_SB_bit_inst_19_n120,
         SD1_SB_inst_SD1_SB_bit_inst_19_n119,
         SD1_SB_inst_SD1_SB_bit_inst_19_n118,
         SD1_SB_inst_SD1_SB_bit_inst_19_n117,
         SD1_SB_inst_SD1_SB_bit_inst_19_n116,
         SD1_SB_inst_SD1_SB_bit_inst_19_n115,
         SD1_SB_inst_SD1_SB_bit_inst_19_n114,
         SD1_SB_inst_SD1_SB_bit_inst_19_n113,
         SD1_SB_inst_SD1_SB_bit_inst_19_n112,
         SD1_SB_inst_SD1_SB_bit_inst_19_n111,
         SD1_SB_inst_SD1_SB_bit_inst_19_n110,
         SD1_SB_inst_SD1_SB_bit_inst_19_n109,
         SD1_SB_inst_SD1_SB_bit_inst_19_n108,
         SD1_SB_inst_SD1_SB_bit_inst_19_n107,
         SD1_SB_inst_SD1_SB_bit_inst_19_n106,
         SD1_SB_inst_SD1_SB_bit_inst_19_n105,
         SD1_SB_inst_SD1_SB_bit_inst_19_n104,
         SD1_SB_inst_SD1_SB_bit_inst_19_n103,
         SD1_SB_inst_SD1_SB_bit_inst_19_n102,
         SD1_SB_inst_SD1_SB_bit_inst_19_n101,
         SD1_SB_inst_SD1_SB_bit_inst_19_n100,
         SD1_SB_inst_SD1_SB_bit_inst_20_n131,
         SD1_SB_inst_SD1_SB_bit_inst_20_n130,
         SD1_SB_inst_SD1_SB_bit_inst_20_n129,
         SD1_SB_inst_SD1_SB_bit_inst_20_n128,
         SD1_SB_inst_SD1_SB_bit_inst_20_n127,
         SD1_SB_inst_SD1_SB_bit_inst_20_n126,
         SD1_SB_inst_SD1_SB_bit_inst_20_n125,
         SD1_SB_inst_SD1_SB_bit_inst_20_n124,
         SD1_SB_inst_SD1_SB_bit_inst_20_n123,
         SD1_SB_inst_SD1_SB_bit_inst_20_n122,
         SD1_SB_inst_SD1_SB_bit_inst_20_n121,
         SD1_SB_inst_SD1_SB_bit_inst_20_n120,
         SD1_SB_inst_SD1_SB_bit_inst_20_n119,
         SD1_SB_inst_SD1_SB_bit_inst_20_n118,
         SD1_SB_inst_SD1_SB_bit_inst_20_n117,
         SD1_SB_inst_SD1_SB_bit_inst_20_n116,
         SD1_SB_inst_SD1_SB_bit_inst_20_n115,
         SD1_SB_inst_SD1_SB_bit_inst_20_n114,
         SD1_SB_inst_SD1_SB_bit_inst_20_n113,
         SD1_SB_inst_SD1_SB_bit_inst_20_n112,
         SD1_SB_inst_SD1_SB_bit_inst_20_n111,
         SD1_SB_inst_SD1_SB_bit_inst_20_n110,
         SD1_SB_inst_SD1_SB_bit_inst_20_n109,
         SD1_SB_inst_SD1_SB_bit_inst_20_n108,
         SD1_SB_inst_SD1_SB_bit_inst_20_n107,
         SD1_SB_inst_SD1_SB_bit_inst_20_n106,
         SD1_SB_inst_SD1_SB_bit_inst_20_n105,
         SD1_SB_inst_SD1_SB_bit_inst_20_n104,
         SD1_SB_inst_SD1_SB_bit_inst_20_n103,
         SD1_SB_inst_SD1_SB_bit_inst_20_n102,
         SD1_SB_inst_SD1_SB_bit_inst_20_n101,
         SD1_SB_inst_SD1_SB_bit_inst_20_n100,
         SD1_SB_inst_SD1_SB_bit_inst_20_n99,
         SD1_SB_inst_SD1_SB_bit_inst_20_n98,
         SD1_SB_inst_SD1_SB_bit_inst_20_n97,
         SD1_SB_inst_SD1_SB_bit_inst_20_n96,
         SD1_SB_inst_SD1_SB_bit_inst_20_n95,
         SD1_SB_inst_SD1_SB_bit_inst_20_n94,
         SD1_SB_inst_SD1_SB_bit_inst_20_n93,
         SD1_SB_inst_SD1_SB_bit_inst_20_n92,
         SD1_SB_inst_SD1_SB_bit_inst_21_n110,
         SD1_SB_inst_SD1_SB_bit_inst_21_n109,
         SD1_SB_inst_SD1_SB_bit_inst_21_n108,
         SD1_SB_inst_SD1_SB_bit_inst_21_n107,
         SD1_SB_inst_SD1_SB_bit_inst_21_n106,
         SD1_SB_inst_SD1_SB_bit_inst_21_n105,
         SD1_SB_inst_SD1_SB_bit_inst_21_n104,
         SD1_SB_inst_SD1_SB_bit_inst_21_n103,
         SD1_SB_inst_SD1_SB_bit_inst_21_n102,
         SD1_SB_inst_SD1_SB_bit_inst_21_n101,
         SD1_SB_inst_SD1_SB_bit_inst_21_n100,
         SD1_SB_inst_SD1_SB_bit_inst_21_n99,
         SD1_SB_inst_SD1_SB_bit_inst_21_n98,
         SD1_SB_inst_SD1_SB_bit_inst_21_n97,
         SD1_SB_inst_SD1_SB_bit_inst_21_n96,
         SD1_SB_inst_SD1_SB_bit_inst_21_n95,
         SD1_SB_inst_SD1_SB_bit_inst_21_n94,
         SD1_SB_inst_SD1_SB_bit_inst_21_n93,
         SD1_SB_inst_SD1_SB_bit_inst_21_n92,
         SD1_SB_inst_SD1_SB_bit_inst_21_n91,
         SD1_SB_inst_SD1_SB_bit_inst_21_n90,
         SD1_SB_inst_SD1_SB_bit_inst_21_n89,
         SD1_SB_inst_SD1_SB_bit_inst_21_n88,
         SD1_SB_inst_SD1_SB_bit_inst_21_n87,
         SD1_SB_inst_SD1_SB_bit_inst_21_n86,
         SD1_SB_inst_SD1_SB_bit_inst_21_n85,
         SD1_SB_inst_SD1_SB_bit_inst_21_n84,
         SD1_SB_inst_SD1_SB_bit_inst_21_n83,
         SD1_SB_inst_SD1_SB_bit_inst_21_n82,
         SD1_SB_inst_SD1_SB_bit_inst_21_n81,
         SD1_SB_inst_SD1_SB_bit_inst_21_n80,
         SD1_SB_inst_SD1_SB_bit_inst_21_n79,
         SD1_SB_inst_SD1_SB_bit_inst_21_n78,
         SD1_SB_inst_SD1_SB_bit_inst_21_n77,
         SD1_SB_inst_SD1_SB_bit_inst_22_n138,
         SD1_SB_inst_SD1_SB_bit_inst_22_n137,
         SD1_SB_inst_SD1_SB_bit_inst_22_n136,
         SD1_SB_inst_SD1_SB_bit_inst_22_n135,
         SD1_SB_inst_SD1_SB_bit_inst_22_n134,
         SD1_SB_inst_SD1_SB_bit_inst_22_n133,
         SD1_SB_inst_SD1_SB_bit_inst_22_n132,
         SD1_SB_inst_SD1_SB_bit_inst_22_n131,
         SD1_SB_inst_SD1_SB_bit_inst_22_n130,
         SD1_SB_inst_SD1_SB_bit_inst_22_n129,
         SD1_SB_inst_SD1_SB_bit_inst_22_n128,
         SD1_SB_inst_SD1_SB_bit_inst_22_n127,
         SD1_SB_inst_SD1_SB_bit_inst_22_n126,
         SD1_SB_inst_SD1_SB_bit_inst_22_n125,
         SD1_SB_inst_SD1_SB_bit_inst_22_n124,
         SD1_SB_inst_SD1_SB_bit_inst_22_n123,
         SD1_SB_inst_SD1_SB_bit_inst_22_n122,
         SD1_SB_inst_SD1_SB_bit_inst_22_n121,
         SD1_SB_inst_SD1_SB_bit_inst_22_n120,
         SD1_SB_inst_SD1_SB_bit_inst_22_n119,
         SD1_SB_inst_SD1_SB_bit_inst_22_n118,
         SD1_SB_inst_SD1_SB_bit_inst_22_n117,
         SD1_SB_inst_SD1_SB_bit_inst_22_n116,
         SD1_SB_inst_SD1_SB_bit_inst_22_n115,
         SD1_SB_inst_SD1_SB_bit_inst_22_n114,
         SD1_SB_inst_SD1_SB_bit_inst_22_n113,
         SD1_SB_inst_SD1_SB_bit_inst_22_n112,
         SD1_SB_inst_SD1_SB_bit_inst_22_n111,
         SD1_SB_inst_SD1_SB_bit_inst_22_n110,
         SD1_SB_inst_SD1_SB_bit_inst_22_n109,
         SD1_SB_inst_SD1_SB_bit_inst_22_n108,
         SD1_SB_inst_SD1_SB_bit_inst_22_n107,
         SD1_SB_inst_SD1_SB_bit_inst_22_n106,
         SD1_SB_inst_SD1_SB_bit_inst_22_n105,
         SD1_SB_inst_SD1_SB_bit_inst_22_n104,
         SD1_SB_inst_SD1_SB_bit_inst_22_n103,
         SD1_SB_inst_SD1_SB_bit_inst_22_n102,
         SD1_SB_inst_SD1_SB_bit_inst_22_n101,
         SD1_SB_inst_SD1_SB_bit_inst_22_n100,
         SD1_SB_inst_SD1_SB_bit_inst_22_n99,
         SD1_SB_inst_SD1_SB_bit_inst_22_n98,
         SD1_SB_inst_SD1_SB_bit_inst_22_n97,
         SD1_SB_inst_SD1_SB_bit_inst_23_n141,
         SD1_SB_inst_SD1_SB_bit_inst_23_n140,
         SD1_SB_inst_SD1_SB_bit_inst_23_n139,
         SD1_SB_inst_SD1_SB_bit_inst_23_n138,
         SD1_SB_inst_SD1_SB_bit_inst_23_n137,
         SD1_SB_inst_SD1_SB_bit_inst_23_n136,
         SD1_SB_inst_SD1_SB_bit_inst_23_n135,
         SD1_SB_inst_SD1_SB_bit_inst_23_n134,
         SD1_SB_inst_SD1_SB_bit_inst_23_n133,
         SD1_SB_inst_SD1_SB_bit_inst_23_n132,
         SD1_SB_inst_SD1_SB_bit_inst_23_n131,
         SD1_SB_inst_SD1_SB_bit_inst_23_n130,
         SD1_SB_inst_SD1_SB_bit_inst_23_n129,
         SD1_SB_inst_SD1_SB_bit_inst_23_n128,
         SD1_SB_inst_SD1_SB_bit_inst_23_n127,
         SD1_SB_inst_SD1_SB_bit_inst_23_n126,
         SD1_SB_inst_SD1_SB_bit_inst_23_n125,
         SD1_SB_inst_SD1_SB_bit_inst_23_n124,
         SD1_SB_inst_SD1_SB_bit_inst_23_n123,
         SD1_SB_inst_SD1_SB_bit_inst_23_n122,
         SD1_SB_inst_SD1_SB_bit_inst_23_n121,
         SD1_SB_inst_SD1_SB_bit_inst_23_n120,
         SD1_SB_inst_SD1_SB_bit_inst_23_n119,
         SD1_SB_inst_SD1_SB_bit_inst_23_n118,
         SD1_SB_inst_SD1_SB_bit_inst_23_n117,
         SD1_SB_inst_SD1_SB_bit_inst_23_n116,
         SD1_SB_inst_SD1_SB_bit_inst_23_n115,
         SD1_SB_inst_SD1_SB_bit_inst_23_n114,
         SD1_SB_inst_SD1_SB_bit_inst_23_n113,
         SD1_SB_inst_SD1_SB_bit_inst_23_n112,
         SD1_SB_inst_SD1_SB_bit_inst_23_n111,
         SD1_SB_inst_SD1_SB_bit_inst_23_n110,
         SD1_SB_inst_SD1_SB_bit_inst_23_n109,
         SD1_SB_inst_SD1_SB_bit_inst_23_n108,
         SD1_SB_inst_SD1_SB_bit_inst_23_n107,
         SD1_SB_inst_SD1_SB_bit_inst_23_n106,
         SD1_SB_inst_SD1_SB_bit_inst_23_n105,
         SD1_SB_inst_SD1_SB_bit_inst_23_n104,
         SD1_SB_inst_SD1_SB_bit_inst_23_n103,
         SD1_SB_inst_SD1_SB_bit_inst_23_n102,
         SD1_SB_inst_SD1_SB_bit_inst_23_n101,
         SD1_SB_inst_SD1_SB_bit_inst_23_n100,
         SD1_SB_inst_SD1_SB_bit_inst_24_n131,
         SD1_SB_inst_SD1_SB_bit_inst_24_n130,
         SD1_SB_inst_SD1_SB_bit_inst_24_n129,
         SD1_SB_inst_SD1_SB_bit_inst_24_n128,
         SD1_SB_inst_SD1_SB_bit_inst_24_n127,
         SD1_SB_inst_SD1_SB_bit_inst_24_n126,
         SD1_SB_inst_SD1_SB_bit_inst_24_n125,
         SD1_SB_inst_SD1_SB_bit_inst_24_n124,
         SD1_SB_inst_SD1_SB_bit_inst_24_n123,
         SD1_SB_inst_SD1_SB_bit_inst_24_n122,
         SD1_SB_inst_SD1_SB_bit_inst_24_n121,
         SD1_SB_inst_SD1_SB_bit_inst_24_n120,
         SD1_SB_inst_SD1_SB_bit_inst_24_n119,
         SD1_SB_inst_SD1_SB_bit_inst_24_n118,
         SD1_SB_inst_SD1_SB_bit_inst_24_n117,
         SD1_SB_inst_SD1_SB_bit_inst_24_n116,
         SD1_SB_inst_SD1_SB_bit_inst_24_n115,
         SD1_SB_inst_SD1_SB_bit_inst_24_n114,
         SD1_SB_inst_SD1_SB_bit_inst_24_n113,
         SD1_SB_inst_SD1_SB_bit_inst_24_n112,
         SD1_SB_inst_SD1_SB_bit_inst_24_n111,
         SD1_SB_inst_SD1_SB_bit_inst_24_n110,
         SD1_SB_inst_SD1_SB_bit_inst_24_n109,
         SD1_SB_inst_SD1_SB_bit_inst_24_n108,
         SD1_SB_inst_SD1_SB_bit_inst_24_n107,
         SD1_SB_inst_SD1_SB_bit_inst_24_n106,
         SD1_SB_inst_SD1_SB_bit_inst_24_n105,
         SD1_SB_inst_SD1_SB_bit_inst_24_n104,
         SD1_SB_inst_SD1_SB_bit_inst_24_n103,
         SD1_SB_inst_SD1_SB_bit_inst_24_n102,
         SD1_SB_inst_SD1_SB_bit_inst_24_n101,
         SD1_SB_inst_SD1_SB_bit_inst_24_n100,
         SD1_SB_inst_SD1_SB_bit_inst_24_n99,
         SD1_SB_inst_SD1_SB_bit_inst_24_n98,
         SD1_SB_inst_SD1_SB_bit_inst_24_n97,
         SD1_SB_inst_SD1_SB_bit_inst_24_n96,
         SD1_SB_inst_SD1_SB_bit_inst_24_n95,
         SD1_SB_inst_SD1_SB_bit_inst_24_n94,
         SD1_SB_inst_SD1_SB_bit_inst_24_n93,
         SD1_SB_inst_SD1_SB_bit_inst_24_n92,
         SD1_SB_inst_SD1_SB_bit_inst_25_n110,
         SD1_SB_inst_SD1_SB_bit_inst_25_n109,
         SD1_SB_inst_SD1_SB_bit_inst_25_n108,
         SD1_SB_inst_SD1_SB_bit_inst_25_n107,
         SD1_SB_inst_SD1_SB_bit_inst_25_n106,
         SD1_SB_inst_SD1_SB_bit_inst_25_n105,
         SD1_SB_inst_SD1_SB_bit_inst_25_n104,
         SD1_SB_inst_SD1_SB_bit_inst_25_n103,
         SD1_SB_inst_SD1_SB_bit_inst_25_n102,
         SD1_SB_inst_SD1_SB_bit_inst_25_n101,
         SD1_SB_inst_SD1_SB_bit_inst_25_n100,
         SD1_SB_inst_SD1_SB_bit_inst_25_n99,
         SD1_SB_inst_SD1_SB_bit_inst_25_n98,
         SD1_SB_inst_SD1_SB_bit_inst_25_n97,
         SD1_SB_inst_SD1_SB_bit_inst_25_n96,
         SD1_SB_inst_SD1_SB_bit_inst_25_n95,
         SD1_SB_inst_SD1_SB_bit_inst_25_n94,
         SD1_SB_inst_SD1_SB_bit_inst_25_n93,
         SD1_SB_inst_SD1_SB_bit_inst_25_n92,
         SD1_SB_inst_SD1_SB_bit_inst_25_n91,
         SD1_SB_inst_SD1_SB_bit_inst_25_n90,
         SD1_SB_inst_SD1_SB_bit_inst_25_n89,
         SD1_SB_inst_SD1_SB_bit_inst_25_n88,
         SD1_SB_inst_SD1_SB_bit_inst_25_n87,
         SD1_SB_inst_SD1_SB_bit_inst_25_n86,
         SD1_SB_inst_SD1_SB_bit_inst_25_n85,
         SD1_SB_inst_SD1_SB_bit_inst_25_n84,
         SD1_SB_inst_SD1_SB_bit_inst_25_n83,
         SD1_SB_inst_SD1_SB_bit_inst_25_n82,
         SD1_SB_inst_SD1_SB_bit_inst_25_n81,
         SD1_SB_inst_SD1_SB_bit_inst_25_n80,
         SD1_SB_inst_SD1_SB_bit_inst_25_n79,
         SD1_SB_inst_SD1_SB_bit_inst_25_n78,
         SD1_SB_inst_SD1_SB_bit_inst_25_n77,
         SD1_SB_inst_SD1_SB_bit_inst_26_n138,
         SD1_SB_inst_SD1_SB_bit_inst_26_n137,
         SD1_SB_inst_SD1_SB_bit_inst_26_n136,
         SD1_SB_inst_SD1_SB_bit_inst_26_n135,
         SD1_SB_inst_SD1_SB_bit_inst_26_n134,
         SD1_SB_inst_SD1_SB_bit_inst_26_n133,
         SD1_SB_inst_SD1_SB_bit_inst_26_n132,
         SD1_SB_inst_SD1_SB_bit_inst_26_n131,
         SD1_SB_inst_SD1_SB_bit_inst_26_n130,
         SD1_SB_inst_SD1_SB_bit_inst_26_n129,
         SD1_SB_inst_SD1_SB_bit_inst_26_n128,
         SD1_SB_inst_SD1_SB_bit_inst_26_n127,
         SD1_SB_inst_SD1_SB_bit_inst_26_n126,
         SD1_SB_inst_SD1_SB_bit_inst_26_n125,
         SD1_SB_inst_SD1_SB_bit_inst_26_n124,
         SD1_SB_inst_SD1_SB_bit_inst_26_n123,
         SD1_SB_inst_SD1_SB_bit_inst_26_n122,
         SD1_SB_inst_SD1_SB_bit_inst_26_n121,
         SD1_SB_inst_SD1_SB_bit_inst_26_n120,
         SD1_SB_inst_SD1_SB_bit_inst_26_n119,
         SD1_SB_inst_SD1_SB_bit_inst_26_n118,
         SD1_SB_inst_SD1_SB_bit_inst_26_n117,
         SD1_SB_inst_SD1_SB_bit_inst_26_n116,
         SD1_SB_inst_SD1_SB_bit_inst_26_n115,
         SD1_SB_inst_SD1_SB_bit_inst_26_n114,
         SD1_SB_inst_SD1_SB_bit_inst_26_n113,
         SD1_SB_inst_SD1_SB_bit_inst_26_n112,
         SD1_SB_inst_SD1_SB_bit_inst_26_n111,
         SD1_SB_inst_SD1_SB_bit_inst_26_n110,
         SD1_SB_inst_SD1_SB_bit_inst_26_n109,
         SD1_SB_inst_SD1_SB_bit_inst_26_n108,
         SD1_SB_inst_SD1_SB_bit_inst_26_n107,
         SD1_SB_inst_SD1_SB_bit_inst_26_n106,
         SD1_SB_inst_SD1_SB_bit_inst_26_n105,
         SD1_SB_inst_SD1_SB_bit_inst_26_n104,
         SD1_SB_inst_SD1_SB_bit_inst_26_n103,
         SD1_SB_inst_SD1_SB_bit_inst_26_n102,
         SD1_SB_inst_SD1_SB_bit_inst_26_n101,
         SD1_SB_inst_SD1_SB_bit_inst_26_n100,
         SD1_SB_inst_SD1_SB_bit_inst_26_n99,
         SD1_SB_inst_SD1_SB_bit_inst_26_n98,
         SD1_SB_inst_SD1_SB_bit_inst_26_n97,
         SD1_SB_inst_SD1_SB_bit_inst_27_n141,
         SD1_SB_inst_SD1_SB_bit_inst_27_n140,
         SD1_SB_inst_SD1_SB_bit_inst_27_n139,
         SD1_SB_inst_SD1_SB_bit_inst_27_n138,
         SD1_SB_inst_SD1_SB_bit_inst_27_n137,
         SD1_SB_inst_SD1_SB_bit_inst_27_n136,
         SD1_SB_inst_SD1_SB_bit_inst_27_n135,
         SD1_SB_inst_SD1_SB_bit_inst_27_n134,
         SD1_SB_inst_SD1_SB_bit_inst_27_n133,
         SD1_SB_inst_SD1_SB_bit_inst_27_n132,
         SD1_SB_inst_SD1_SB_bit_inst_27_n131,
         SD1_SB_inst_SD1_SB_bit_inst_27_n130,
         SD1_SB_inst_SD1_SB_bit_inst_27_n129,
         SD1_SB_inst_SD1_SB_bit_inst_27_n128,
         SD1_SB_inst_SD1_SB_bit_inst_27_n127,
         SD1_SB_inst_SD1_SB_bit_inst_27_n126,
         SD1_SB_inst_SD1_SB_bit_inst_27_n125,
         SD1_SB_inst_SD1_SB_bit_inst_27_n124,
         SD1_SB_inst_SD1_SB_bit_inst_27_n123,
         SD1_SB_inst_SD1_SB_bit_inst_27_n122,
         SD1_SB_inst_SD1_SB_bit_inst_27_n121,
         SD1_SB_inst_SD1_SB_bit_inst_27_n120,
         SD1_SB_inst_SD1_SB_bit_inst_27_n119,
         SD1_SB_inst_SD1_SB_bit_inst_27_n118,
         SD1_SB_inst_SD1_SB_bit_inst_27_n117,
         SD1_SB_inst_SD1_SB_bit_inst_27_n116,
         SD1_SB_inst_SD1_SB_bit_inst_27_n115,
         SD1_SB_inst_SD1_SB_bit_inst_27_n114,
         SD1_SB_inst_SD1_SB_bit_inst_27_n113,
         SD1_SB_inst_SD1_SB_bit_inst_27_n112,
         SD1_SB_inst_SD1_SB_bit_inst_27_n111,
         SD1_SB_inst_SD1_SB_bit_inst_27_n110,
         SD1_SB_inst_SD1_SB_bit_inst_27_n109,
         SD1_SB_inst_SD1_SB_bit_inst_27_n108,
         SD1_SB_inst_SD1_SB_bit_inst_27_n107,
         SD1_SB_inst_SD1_SB_bit_inst_27_n106,
         SD1_SB_inst_SD1_SB_bit_inst_27_n105,
         SD1_SB_inst_SD1_SB_bit_inst_27_n104,
         SD1_SB_inst_SD1_SB_bit_inst_27_n103,
         SD1_SB_inst_SD1_SB_bit_inst_27_n102,
         SD1_SB_inst_SD1_SB_bit_inst_27_n101,
         SD1_SB_inst_SD1_SB_bit_inst_27_n100,
         SD1_SB_inst_SD1_SB_bit_inst_28_n132,
         SD1_SB_inst_SD1_SB_bit_inst_28_n131,
         SD1_SB_inst_SD1_SB_bit_inst_28_n130,
         SD1_SB_inst_SD1_SB_bit_inst_28_n129,
         SD1_SB_inst_SD1_SB_bit_inst_28_n128,
         SD1_SB_inst_SD1_SB_bit_inst_28_n127,
         SD1_SB_inst_SD1_SB_bit_inst_28_n126,
         SD1_SB_inst_SD1_SB_bit_inst_28_n125,
         SD1_SB_inst_SD1_SB_bit_inst_28_n124,
         SD1_SB_inst_SD1_SB_bit_inst_28_n123,
         SD1_SB_inst_SD1_SB_bit_inst_28_n122,
         SD1_SB_inst_SD1_SB_bit_inst_28_n121,
         SD1_SB_inst_SD1_SB_bit_inst_28_n120,
         SD1_SB_inst_SD1_SB_bit_inst_28_n119,
         SD1_SB_inst_SD1_SB_bit_inst_28_n118,
         SD1_SB_inst_SD1_SB_bit_inst_28_n117,
         SD1_SB_inst_SD1_SB_bit_inst_28_n116,
         SD1_SB_inst_SD1_SB_bit_inst_28_n115,
         SD1_SB_inst_SD1_SB_bit_inst_28_n114,
         SD1_SB_inst_SD1_SB_bit_inst_28_n113,
         SD1_SB_inst_SD1_SB_bit_inst_28_n112,
         SD1_SB_inst_SD1_SB_bit_inst_28_n111,
         SD1_SB_inst_SD1_SB_bit_inst_28_n110,
         SD1_SB_inst_SD1_SB_bit_inst_28_n109,
         SD1_SB_inst_SD1_SB_bit_inst_28_n108,
         SD1_SB_inst_SD1_SB_bit_inst_28_n107,
         SD1_SB_inst_SD1_SB_bit_inst_28_n106,
         SD1_SB_inst_SD1_SB_bit_inst_28_n105,
         SD1_SB_inst_SD1_SB_bit_inst_28_n104,
         SD1_SB_inst_SD1_SB_bit_inst_28_n103,
         SD1_SB_inst_SD1_SB_bit_inst_28_n102,
         SD1_SB_inst_SD1_SB_bit_inst_28_n101,
         SD1_SB_inst_SD1_SB_bit_inst_28_n100,
         SD1_SB_inst_SD1_SB_bit_inst_28_n99,
         SD1_SB_inst_SD1_SB_bit_inst_28_n98,
         SD1_SB_inst_SD1_SB_bit_inst_28_n97,
         SD1_SB_inst_SD1_SB_bit_inst_28_n96,
         SD1_SB_inst_SD1_SB_bit_inst_28_n95,
         SD1_SB_inst_SD1_SB_bit_inst_28_n94,
         SD1_SB_inst_SD1_SB_bit_inst_28_n93,
         SD1_SB_inst_SD1_SB_bit_inst_28_n92,
         SD1_SB_inst_SD1_SB_bit_inst_29_n109,
         SD1_SB_inst_SD1_SB_bit_inst_29_n108,
         SD1_SB_inst_SD1_SB_bit_inst_29_n107,
         SD1_SB_inst_SD1_SB_bit_inst_29_n106,
         SD1_SB_inst_SD1_SB_bit_inst_29_n105,
         SD1_SB_inst_SD1_SB_bit_inst_29_n104,
         SD1_SB_inst_SD1_SB_bit_inst_29_n103,
         SD1_SB_inst_SD1_SB_bit_inst_29_n102,
         SD1_SB_inst_SD1_SB_bit_inst_29_n101,
         SD1_SB_inst_SD1_SB_bit_inst_29_n100,
         SD1_SB_inst_SD1_SB_bit_inst_29_n99,
         SD1_SB_inst_SD1_SB_bit_inst_29_n98,
         SD1_SB_inst_SD1_SB_bit_inst_29_n97,
         SD1_SB_inst_SD1_SB_bit_inst_29_n96,
         SD1_SB_inst_SD1_SB_bit_inst_29_n95,
         SD1_SB_inst_SD1_SB_bit_inst_29_n94,
         SD1_SB_inst_SD1_SB_bit_inst_29_n93,
         SD1_SB_inst_SD1_SB_bit_inst_29_n92,
         SD1_SB_inst_SD1_SB_bit_inst_29_n91,
         SD1_SB_inst_SD1_SB_bit_inst_29_n90,
         SD1_SB_inst_SD1_SB_bit_inst_29_n89,
         SD1_SB_inst_SD1_SB_bit_inst_29_n88,
         SD1_SB_inst_SD1_SB_bit_inst_29_n87,
         SD1_SB_inst_SD1_SB_bit_inst_29_n86,
         SD1_SB_inst_SD1_SB_bit_inst_29_n85,
         SD1_SB_inst_SD1_SB_bit_inst_29_n84,
         SD1_SB_inst_SD1_SB_bit_inst_29_n83,
         SD1_SB_inst_SD1_SB_bit_inst_29_n82,
         SD1_SB_inst_SD1_SB_bit_inst_29_n81,
         SD1_SB_inst_SD1_SB_bit_inst_29_n80,
         SD1_SB_inst_SD1_SB_bit_inst_29_n79,
         SD1_SB_inst_SD1_SB_bit_inst_29_n78,
         SD1_SB_inst_SD1_SB_bit_inst_29_n77,
         SD1_SB_inst_SD1_SB_bit_inst_30_n137,
         SD1_SB_inst_SD1_SB_bit_inst_30_n136,
         SD1_SB_inst_SD1_SB_bit_inst_30_n135,
         SD1_SB_inst_SD1_SB_bit_inst_30_n134,
         SD1_SB_inst_SD1_SB_bit_inst_30_n133,
         SD1_SB_inst_SD1_SB_bit_inst_30_n132,
         SD1_SB_inst_SD1_SB_bit_inst_30_n131,
         SD1_SB_inst_SD1_SB_bit_inst_30_n130,
         SD1_SB_inst_SD1_SB_bit_inst_30_n129,
         SD1_SB_inst_SD1_SB_bit_inst_30_n128,
         SD1_SB_inst_SD1_SB_bit_inst_30_n127,
         SD1_SB_inst_SD1_SB_bit_inst_30_n126,
         SD1_SB_inst_SD1_SB_bit_inst_30_n125,
         SD1_SB_inst_SD1_SB_bit_inst_30_n124,
         SD1_SB_inst_SD1_SB_bit_inst_30_n123,
         SD1_SB_inst_SD1_SB_bit_inst_30_n122,
         SD1_SB_inst_SD1_SB_bit_inst_30_n121,
         SD1_SB_inst_SD1_SB_bit_inst_30_n120,
         SD1_SB_inst_SD1_SB_bit_inst_30_n119,
         SD1_SB_inst_SD1_SB_bit_inst_30_n118,
         SD1_SB_inst_SD1_SB_bit_inst_30_n117,
         SD1_SB_inst_SD1_SB_bit_inst_30_n116,
         SD1_SB_inst_SD1_SB_bit_inst_30_n115,
         SD1_SB_inst_SD1_SB_bit_inst_30_n114,
         SD1_SB_inst_SD1_SB_bit_inst_30_n113,
         SD1_SB_inst_SD1_SB_bit_inst_30_n112,
         SD1_SB_inst_SD1_SB_bit_inst_30_n111,
         SD1_SB_inst_SD1_SB_bit_inst_30_n110,
         SD1_SB_inst_SD1_SB_bit_inst_30_n109,
         SD1_SB_inst_SD1_SB_bit_inst_30_n108,
         SD1_SB_inst_SD1_SB_bit_inst_30_n107,
         SD1_SB_inst_SD1_SB_bit_inst_30_n106,
         SD1_SB_inst_SD1_SB_bit_inst_30_n105,
         SD1_SB_inst_SD1_SB_bit_inst_30_n104,
         SD1_SB_inst_SD1_SB_bit_inst_30_n103,
         SD1_SB_inst_SD1_SB_bit_inst_30_n102,
         SD1_SB_inst_SD1_SB_bit_inst_30_n101,
         SD1_SB_inst_SD1_SB_bit_inst_30_n100,
         SD1_SB_inst_SD1_SB_bit_inst_30_n99,
         SD1_SB_inst_SD1_SB_bit_inst_30_n98,
         SD1_SB_inst_SD1_SB_bit_inst_30_n97,
         SD1_SB_inst_SD1_SB_bit_inst_31_n141,
         SD1_SB_inst_SD1_SB_bit_inst_31_n140,
         SD1_SB_inst_SD1_SB_bit_inst_31_n139,
         SD1_SB_inst_SD1_SB_bit_inst_31_n138,
         SD1_SB_inst_SD1_SB_bit_inst_31_n137,
         SD1_SB_inst_SD1_SB_bit_inst_31_n136,
         SD1_SB_inst_SD1_SB_bit_inst_31_n135,
         SD1_SB_inst_SD1_SB_bit_inst_31_n134,
         SD1_SB_inst_SD1_SB_bit_inst_31_n133,
         SD1_SB_inst_SD1_SB_bit_inst_31_n132,
         SD1_SB_inst_SD1_SB_bit_inst_31_n131,
         SD1_SB_inst_SD1_SB_bit_inst_31_n130,
         SD1_SB_inst_SD1_SB_bit_inst_31_n129,
         SD1_SB_inst_SD1_SB_bit_inst_31_n128,
         SD1_SB_inst_SD1_SB_bit_inst_31_n127,
         SD1_SB_inst_SD1_SB_bit_inst_31_n126,
         SD1_SB_inst_SD1_SB_bit_inst_31_n125,
         SD1_SB_inst_SD1_SB_bit_inst_31_n124,
         SD1_SB_inst_SD1_SB_bit_inst_31_n123,
         SD1_SB_inst_SD1_SB_bit_inst_31_n122,
         SD1_SB_inst_SD1_SB_bit_inst_31_n121,
         SD1_SB_inst_SD1_SB_bit_inst_31_n120,
         SD1_SB_inst_SD1_SB_bit_inst_31_n119,
         SD1_SB_inst_SD1_SB_bit_inst_31_n118,
         SD1_SB_inst_SD1_SB_bit_inst_31_n117,
         SD1_SB_inst_SD1_SB_bit_inst_31_n116,
         SD1_SB_inst_SD1_SB_bit_inst_31_n115,
         SD1_SB_inst_SD1_SB_bit_inst_31_n114,
         SD1_SB_inst_SD1_SB_bit_inst_31_n113,
         SD1_SB_inst_SD1_SB_bit_inst_31_n112,
         SD1_SB_inst_SD1_SB_bit_inst_31_n111,
         SD1_SB_inst_SD1_SB_bit_inst_31_n110,
         SD1_SB_inst_SD1_SB_bit_inst_31_n109,
         SD1_SB_inst_SD1_SB_bit_inst_31_n108,
         SD1_SB_inst_SD1_SB_bit_inst_31_n107,
         SD1_SB_inst_SD1_SB_bit_inst_31_n106,
         SD1_SB_inst_SD1_SB_bit_inst_31_n105,
         SD1_SB_inst_SD1_SB_bit_inst_31_n104,
         SD1_SB_inst_SD1_SB_bit_inst_31_n103,
         SD1_SB_inst_SD1_SB_bit_inst_31_n102,
         SD1_SB_inst_SD1_SB_bit_inst_31_n101,
         SD1_SB_inst_SD1_SB_bit_inst_31_n100,
         SD1_SB_inst_SD1_SB_bit_inst_32_n131,
         SD1_SB_inst_SD1_SB_bit_inst_32_n130,
         SD1_SB_inst_SD1_SB_bit_inst_32_n129,
         SD1_SB_inst_SD1_SB_bit_inst_32_n128,
         SD1_SB_inst_SD1_SB_bit_inst_32_n127,
         SD1_SB_inst_SD1_SB_bit_inst_32_n126,
         SD1_SB_inst_SD1_SB_bit_inst_32_n125,
         SD1_SB_inst_SD1_SB_bit_inst_32_n124,
         SD1_SB_inst_SD1_SB_bit_inst_32_n123,
         SD1_SB_inst_SD1_SB_bit_inst_32_n122,
         SD1_SB_inst_SD1_SB_bit_inst_32_n121,
         SD1_SB_inst_SD1_SB_bit_inst_32_n120,
         SD1_SB_inst_SD1_SB_bit_inst_32_n119,
         SD1_SB_inst_SD1_SB_bit_inst_32_n118,
         SD1_SB_inst_SD1_SB_bit_inst_32_n117,
         SD1_SB_inst_SD1_SB_bit_inst_32_n116,
         SD1_SB_inst_SD1_SB_bit_inst_32_n115,
         SD1_SB_inst_SD1_SB_bit_inst_32_n114,
         SD1_SB_inst_SD1_SB_bit_inst_32_n113,
         SD1_SB_inst_SD1_SB_bit_inst_32_n112,
         SD1_SB_inst_SD1_SB_bit_inst_32_n111,
         SD1_SB_inst_SD1_SB_bit_inst_32_n110,
         SD1_SB_inst_SD1_SB_bit_inst_32_n109,
         SD1_SB_inst_SD1_SB_bit_inst_32_n108,
         SD1_SB_inst_SD1_SB_bit_inst_32_n107,
         SD1_SB_inst_SD1_SB_bit_inst_32_n106,
         SD1_SB_inst_SD1_SB_bit_inst_32_n105,
         SD1_SB_inst_SD1_SB_bit_inst_32_n104,
         SD1_SB_inst_SD1_SB_bit_inst_32_n103,
         SD1_SB_inst_SD1_SB_bit_inst_32_n102,
         SD1_SB_inst_SD1_SB_bit_inst_32_n101,
         SD1_SB_inst_SD1_SB_bit_inst_32_n100,
         SD1_SB_inst_SD1_SB_bit_inst_32_n99,
         SD1_SB_inst_SD1_SB_bit_inst_32_n98,
         SD1_SB_inst_SD1_SB_bit_inst_32_n97,
         SD1_SB_inst_SD1_SB_bit_inst_32_n96,
         SD1_SB_inst_SD1_SB_bit_inst_32_n95,
         SD1_SB_inst_SD1_SB_bit_inst_32_n94,
         SD1_SB_inst_SD1_SB_bit_inst_32_n93,
         SD1_SB_inst_SD1_SB_bit_inst_32_n92,
         SD1_SB_inst_SD1_SB_bit_inst_33_n110,
         SD1_SB_inst_SD1_SB_bit_inst_33_n109,
         SD1_SB_inst_SD1_SB_bit_inst_33_n108,
         SD1_SB_inst_SD1_SB_bit_inst_33_n107,
         SD1_SB_inst_SD1_SB_bit_inst_33_n106,
         SD1_SB_inst_SD1_SB_bit_inst_33_n105,
         SD1_SB_inst_SD1_SB_bit_inst_33_n104,
         SD1_SB_inst_SD1_SB_bit_inst_33_n103,
         SD1_SB_inst_SD1_SB_bit_inst_33_n102,
         SD1_SB_inst_SD1_SB_bit_inst_33_n101,
         SD1_SB_inst_SD1_SB_bit_inst_33_n100,
         SD1_SB_inst_SD1_SB_bit_inst_33_n99,
         SD1_SB_inst_SD1_SB_bit_inst_33_n98,
         SD1_SB_inst_SD1_SB_bit_inst_33_n97,
         SD1_SB_inst_SD1_SB_bit_inst_33_n96,
         SD1_SB_inst_SD1_SB_bit_inst_33_n95,
         SD1_SB_inst_SD1_SB_bit_inst_33_n94,
         SD1_SB_inst_SD1_SB_bit_inst_33_n93,
         SD1_SB_inst_SD1_SB_bit_inst_33_n92,
         SD1_SB_inst_SD1_SB_bit_inst_33_n91,
         SD1_SB_inst_SD1_SB_bit_inst_33_n90,
         SD1_SB_inst_SD1_SB_bit_inst_33_n89,
         SD1_SB_inst_SD1_SB_bit_inst_33_n88,
         SD1_SB_inst_SD1_SB_bit_inst_33_n87,
         SD1_SB_inst_SD1_SB_bit_inst_33_n86,
         SD1_SB_inst_SD1_SB_bit_inst_33_n85,
         SD1_SB_inst_SD1_SB_bit_inst_33_n84,
         SD1_SB_inst_SD1_SB_bit_inst_33_n83,
         SD1_SB_inst_SD1_SB_bit_inst_33_n82,
         SD1_SB_inst_SD1_SB_bit_inst_33_n81,
         SD1_SB_inst_SD1_SB_bit_inst_33_n80,
         SD1_SB_inst_SD1_SB_bit_inst_33_n79,
         SD1_SB_inst_SD1_SB_bit_inst_33_n78,
         SD1_SB_inst_SD1_SB_bit_inst_33_n77,
         SD1_SB_inst_SD1_SB_bit_inst_34_n138,
         SD1_SB_inst_SD1_SB_bit_inst_34_n137,
         SD1_SB_inst_SD1_SB_bit_inst_34_n136,
         SD1_SB_inst_SD1_SB_bit_inst_34_n135,
         SD1_SB_inst_SD1_SB_bit_inst_34_n134,
         SD1_SB_inst_SD1_SB_bit_inst_34_n133,
         SD1_SB_inst_SD1_SB_bit_inst_34_n132,
         SD1_SB_inst_SD1_SB_bit_inst_34_n131,
         SD1_SB_inst_SD1_SB_bit_inst_34_n130,
         SD1_SB_inst_SD1_SB_bit_inst_34_n129,
         SD1_SB_inst_SD1_SB_bit_inst_34_n128,
         SD1_SB_inst_SD1_SB_bit_inst_34_n127,
         SD1_SB_inst_SD1_SB_bit_inst_34_n126,
         SD1_SB_inst_SD1_SB_bit_inst_34_n125,
         SD1_SB_inst_SD1_SB_bit_inst_34_n124,
         SD1_SB_inst_SD1_SB_bit_inst_34_n123,
         SD1_SB_inst_SD1_SB_bit_inst_34_n122,
         SD1_SB_inst_SD1_SB_bit_inst_34_n121,
         SD1_SB_inst_SD1_SB_bit_inst_34_n120,
         SD1_SB_inst_SD1_SB_bit_inst_34_n119,
         SD1_SB_inst_SD1_SB_bit_inst_34_n118,
         SD1_SB_inst_SD1_SB_bit_inst_34_n117,
         SD1_SB_inst_SD1_SB_bit_inst_34_n116,
         SD1_SB_inst_SD1_SB_bit_inst_34_n115,
         SD1_SB_inst_SD1_SB_bit_inst_34_n114,
         SD1_SB_inst_SD1_SB_bit_inst_34_n113,
         SD1_SB_inst_SD1_SB_bit_inst_34_n112,
         SD1_SB_inst_SD1_SB_bit_inst_34_n111,
         SD1_SB_inst_SD1_SB_bit_inst_34_n110,
         SD1_SB_inst_SD1_SB_bit_inst_34_n109,
         SD1_SB_inst_SD1_SB_bit_inst_34_n108,
         SD1_SB_inst_SD1_SB_bit_inst_34_n107,
         SD1_SB_inst_SD1_SB_bit_inst_34_n106,
         SD1_SB_inst_SD1_SB_bit_inst_34_n105,
         SD1_SB_inst_SD1_SB_bit_inst_34_n104,
         SD1_SB_inst_SD1_SB_bit_inst_34_n103,
         SD1_SB_inst_SD1_SB_bit_inst_34_n102,
         SD1_SB_inst_SD1_SB_bit_inst_34_n101,
         SD1_SB_inst_SD1_SB_bit_inst_34_n100,
         SD1_SB_inst_SD1_SB_bit_inst_34_n99,
         SD1_SB_inst_SD1_SB_bit_inst_34_n98,
         SD1_SB_inst_SD1_SB_bit_inst_34_n97,
         SD1_SB_inst_SD1_SB_bit_inst_35_n141,
         SD1_SB_inst_SD1_SB_bit_inst_35_n140,
         SD1_SB_inst_SD1_SB_bit_inst_35_n139,
         SD1_SB_inst_SD1_SB_bit_inst_35_n138,
         SD1_SB_inst_SD1_SB_bit_inst_35_n137,
         SD1_SB_inst_SD1_SB_bit_inst_35_n136,
         SD1_SB_inst_SD1_SB_bit_inst_35_n135,
         SD1_SB_inst_SD1_SB_bit_inst_35_n134,
         SD1_SB_inst_SD1_SB_bit_inst_35_n133,
         SD1_SB_inst_SD1_SB_bit_inst_35_n132,
         SD1_SB_inst_SD1_SB_bit_inst_35_n131,
         SD1_SB_inst_SD1_SB_bit_inst_35_n130,
         SD1_SB_inst_SD1_SB_bit_inst_35_n129,
         SD1_SB_inst_SD1_SB_bit_inst_35_n128,
         SD1_SB_inst_SD1_SB_bit_inst_35_n127,
         SD1_SB_inst_SD1_SB_bit_inst_35_n126,
         SD1_SB_inst_SD1_SB_bit_inst_35_n125,
         SD1_SB_inst_SD1_SB_bit_inst_35_n124,
         SD1_SB_inst_SD1_SB_bit_inst_35_n123,
         SD1_SB_inst_SD1_SB_bit_inst_35_n122,
         SD1_SB_inst_SD1_SB_bit_inst_35_n121,
         SD1_SB_inst_SD1_SB_bit_inst_35_n120,
         SD1_SB_inst_SD1_SB_bit_inst_35_n119,
         SD1_SB_inst_SD1_SB_bit_inst_35_n118,
         SD1_SB_inst_SD1_SB_bit_inst_35_n117,
         SD1_SB_inst_SD1_SB_bit_inst_35_n116,
         SD1_SB_inst_SD1_SB_bit_inst_35_n115,
         SD1_SB_inst_SD1_SB_bit_inst_35_n114,
         SD1_SB_inst_SD1_SB_bit_inst_35_n113,
         SD1_SB_inst_SD1_SB_bit_inst_35_n112,
         SD1_SB_inst_SD1_SB_bit_inst_35_n111,
         SD1_SB_inst_SD1_SB_bit_inst_35_n110,
         SD1_SB_inst_SD1_SB_bit_inst_35_n109,
         SD1_SB_inst_SD1_SB_bit_inst_35_n108,
         SD1_SB_inst_SD1_SB_bit_inst_35_n107,
         SD1_SB_inst_SD1_SB_bit_inst_35_n106,
         SD1_SB_inst_SD1_SB_bit_inst_35_n105,
         SD1_SB_inst_SD1_SB_bit_inst_35_n104,
         SD1_SB_inst_SD1_SB_bit_inst_35_n103,
         SD1_SB_inst_SD1_SB_bit_inst_35_n102,
         SD1_SB_inst_SD1_SB_bit_inst_35_n101,
         SD1_SB_inst_SD1_SB_bit_inst_35_n100,
         SD1_SB_inst_SD1_SB_bit_inst_36_n131,
         SD1_SB_inst_SD1_SB_bit_inst_36_n130,
         SD1_SB_inst_SD1_SB_bit_inst_36_n129,
         SD1_SB_inst_SD1_SB_bit_inst_36_n128,
         SD1_SB_inst_SD1_SB_bit_inst_36_n127,
         SD1_SB_inst_SD1_SB_bit_inst_36_n126,
         SD1_SB_inst_SD1_SB_bit_inst_36_n125,
         SD1_SB_inst_SD1_SB_bit_inst_36_n124,
         SD1_SB_inst_SD1_SB_bit_inst_36_n123,
         SD1_SB_inst_SD1_SB_bit_inst_36_n122,
         SD1_SB_inst_SD1_SB_bit_inst_36_n121,
         SD1_SB_inst_SD1_SB_bit_inst_36_n120,
         SD1_SB_inst_SD1_SB_bit_inst_36_n119,
         SD1_SB_inst_SD1_SB_bit_inst_36_n118,
         SD1_SB_inst_SD1_SB_bit_inst_36_n117,
         SD1_SB_inst_SD1_SB_bit_inst_36_n116,
         SD1_SB_inst_SD1_SB_bit_inst_36_n115,
         SD1_SB_inst_SD1_SB_bit_inst_36_n114,
         SD1_SB_inst_SD1_SB_bit_inst_36_n113,
         SD1_SB_inst_SD1_SB_bit_inst_36_n112,
         SD1_SB_inst_SD1_SB_bit_inst_36_n111,
         SD1_SB_inst_SD1_SB_bit_inst_36_n110,
         SD1_SB_inst_SD1_SB_bit_inst_36_n109,
         SD1_SB_inst_SD1_SB_bit_inst_36_n108,
         SD1_SB_inst_SD1_SB_bit_inst_36_n107,
         SD1_SB_inst_SD1_SB_bit_inst_36_n106,
         SD1_SB_inst_SD1_SB_bit_inst_36_n105,
         SD1_SB_inst_SD1_SB_bit_inst_36_n104,
         SD1_SB_inst_SD1_SB_bit_inst_36_n103,
         SD1_SB_inst_SD1_SB_bit_inst_36_n102,
         SD1_SB_inst_SD1_SB_bit_inst_36_n101,
         SD1_SB_inst_SD1_SB_bit_inst_36_n100,
         SD1_SB_inst_SD1_SB_bit_inst_36_n99,
         SD1_SB_inst_SD1_SB_bit_inst_36_n98,
         SD1_SB_inst_SD1_SB_bit_inst_36_n97,
         SD1_SB_inst_SD1_SB_bit_inst_36_n96,
         SD1_SB_inst_SD1_SB_bit_inst_36_n95,
         SD1_SB_inst_SD1_SB_bit_inst_36_n94,
         SD1_SB_inst_SD1_SB_bit_inst_36_n93,
         SD1_SB_inst_SD1_SB_bit_inst_36_n92,
         SD1_SB_inst_SD1_SB_bit_inst_37_n110,
         SD1_SB_inst_SD1_SB_bit_inst_37_n109,
         SD1_SB_inst_SD1_SB_bit_inst_37_n108,
         SD1_SB_inst_SD1_SB_bit_inst_37_n107,
         SD1_SB_inst_SD1_SB_bit_inst_37_n106,
         SD1_SB_inst_SD1_SB_bit_inst_37_n105,
         SD1_SB_inst_SD1_SB_bit_inst_37_n104,
         SD1_SB_inst_SD1_SB_bit_inst_37_n103,
         SD1_SB_inst_SD1_SB_bit_inst_37_n102,
         SD1_SB_inst_SD1_SB_bit_inst_37_n101,
         SD1_SB_inst_SD1_SB_bit_inst_37_n100,
         SD1_SB_inst_SD1_SB_bit_inst_37_n99,
         SD1_SB_inst_SD1_SB_bit_inst_37_n98,
         SD1_SB_inst_SD1_SB_bit_inst_37_n97,
         SD1_SB_inst_SD1_SB_bit_inst_37_n96,
         SD1_SB_inst_SD1_SB_bit_inst_37_n95,
         SD1_SB_inst_SD1_SB_bit_inst_37_n94,
         SD1_SB_inst_SD1_SB_bit_inst_37_n93,
         SD1_SB_inst_SD1_SB_bit_inst_37_n92,
         SD1_SB_inst_SD1_SB_bit_inst_37_n91,
         SD1_SB_inst_SD1_SB_bit_inst_37_n90,
         SD1_SB_inst_SD1_SB_bit_inst_37_n89,
         SD1_SB_inst_SD1_SB_bit_inst_37_n88,
         SD1_SB_inst_SD1_SB_bit_inst_37_n87,
         SD1_SB_inst_SD1_SB_bit_inst_37_n86,
         SD1_SB_inst_SD1_SB_bit_inst_37_n85,
         SD1_SB_inst_SD1_SB_bit_inst_37_n84,
         SD1_SB_inst_SD1_SB_bit_inst_37_n83,
         SD1_SB_inst_SD1_SB_bit_inst_37_n82,
         SD1_SB_inst_SD1_SB_bit_inst_37_n81,
         SD1_SB_inst_SD1_SB_bit_inst_37_n80,
         SD1_SB_inst_SD1_SB_bit_inst_37_n79,
         SD1_SB_inst_SD1_SB_bit_inst_37_n78,
         SD1_SB_inst_SD1_SB_bit_inst_37_n77,
         SD1_SB_inst_SD1_SB_bit_inst_38_n138,
         SD1_SB_inst_SD1_SB_bit_inst_38_n137,
         SD1_SB_inst_SD1_SB_bit_inst_38_n136,
         SD1_SB_inst_SD1_SB_bit_inst_38_n135,
         SD1_SB_inst_SD1_SB_bit_inst_38_n134,
         SD1_SB_inst_SD1_SB_bit_inst_38_n133,
         SD1_SB_inst_SD1_SB_bit_inst_38_n132,
         SD1_SB_inst_SD1_SB_bit_inst_38_n131,
         SD1_SB_inst_SD1_SB_bit_inst_38_n130,
         SD1_SB_inst_SD1_SB_bit_inst_38_n129,
         SD1_SB_inst_SD1_SB_bit_inst_38_n128,
         SD1_SB_inst_SD1_SB_bit_inst_38_n127,
         SD1_SB_inst_SD1_SB_bit_inst_38_n126,
         SD1_SB_inst_SD1_SB_bit_inst_38_n125,
         SD1_SB_inst_SD1_SB_bit_inst_38_n124,
         SD1_SB_inst_SD1_SB_bit_inst_38_n123,
         SD1_SB_inst_SD1_SB_bit_inst_38_n122,
         SD1_SB_inst_SD1_SB_bit_inst_38_n121,
         SD1_SB_inst_SD1_SB_bit_inst_38_n120,
         SD1_SB_inst_SD1_SB_bit_inst_38_n119,
         SD1_SB_inst_SD1_SB_bit_inst_38_n118,
         SD1_SB_inst_SD1_SB_bit_inst_38_n117,
         SD1_SB_inst_SD1_SB_bit_inst_38_n116,
         SD1_SB_inst_SD1_SB_bit_inst_38_n115,
         SD1_SB_inst_SD1_SB_bit_inst_38_n114,
         SD1_SB_inst_SD1_SB_bit_inst_38_n113,
         SD1_SB_inst_SD1_SB_bit_inst_38_n112,
         SD1_SB_inst_SD1_SB_bit_inst_38_n111,
         SD1_SB_inst_SD1_SB_bit_inst_38_n110,
         SD1_SB_inst_SD1_SB_bit_inst_38_n109,
         SD1_SB_inst_SD1_SB_bit_inst_38_n108,
         SD1_SB_inst_SD1_SB_bit_inst_38_n107,
         SD1_SB_inst_SD1_SB_bit_inst_38_n106,
         SD1_SB_inst_SD1_SB_bit_inst_38_n105,
         SD1_SB_inst_SD1_SB_bit_inst_38_n104,
         SD1_SB_inst_SD1_SB_bit_inst_38_n103,
         SD1_SB_inst_SD1_SB_bit_inst_38_n102,
         SD1_SB_inst_SD1_SB_bit_inst_38_n101,
         SD1_SB_inst_SD1_SB_bit_inst_38_n100,
         SD1_SB_inst_SD1_SB_bit_inst_38_n99,
         SD1_SB_inst_SD1_SB_bit_inst_38_n98,
         SD1_SB_inst_SD1_SB_bit_inst_38_n97,
         SD1_SB_inst_SD1_SB_bit_inst_39_n141,
         SD1_SB_inst_SD1_SB_bit_inst_39_n140,
         SD1_SB_inst_SD1_SB_bit_inst_39_n139,
         SD1_SB_inst_SD1_SB_bit_inst_39_n138,
         SD1_SB_inst_SD1_SB_bit_inst_39_n137,
         SD1_SB_inst_SD1_SB_bit_inst_39_n136,
         SD1_SB_inst_SD1_SB_bit_inst_39_n135,
         SD1_SB_inst_SD1_SB_bit_inst_39_n134,
         SD1_SB_inst_SD1_SB_bit_inst_39_n133,
         SD1_SB_inst_SD1_SB_bit_inst_39_n132,
         SD1_SB_inst_SD1_SB_bit_inst_39_n131,
         SD1_SB_inst_SD1_SB_bit_inst_39_n130,
         SD1_SB_inst_SD1_SB_bit_inst_39_n129,
         SD1_SB_inst_SD1_SB_bit_inst_39_n128,
         SD1_SB_inst_SD1_SB_bit_inst_39_n127,
         SD1_SB_inst_SD1_SB_bit_inst_39_n126,
         SD1_SB_inst_SD1_SB_bit_inst_39_n125,
         SD1_SB_inst_SD1_SB_bit_inst_39_n124,
         SD1_SB_inst_SD1_SB_bit_inst_39_n123,
         SD1_SB_inst_SD1_SB_bit_inst_39_n122,
         SD1_SB_inst_SD1_SB_bit_inst_39_n121,
         SD1_SB_inst_SD1_SB_bit_inst_39_n120,
         SD1_SB_inst_SD1_SB_bit_inst_39_n119,
         SD1_SB_inst_SD1_SB_bit_inst_39_n118,
         SD1_SB_inst_SD1_SB_bit_inst_39_n117,
         SD1_SB_inst_SD1_SB_bit_inst_39_n116,
         SD1_SB_inst_SD1_SB_bit_inst_39_n115,
         SD1_SB_inst_SD1_SB_bit_inst_39_n114,
         SD1_SB_inst_SD1_SB_bit_inst_39_n113,
         SD1_SB_inst_SD1_SB_bit_inst_39_n112,
         SD1_SB_inst_SD1_SB_bit_inst_39_n111,
         SD1_SB_inst_SD1_SB_bit_inst_39_n110,
         SD1_SB_inst_SD1_SB_bit_inst_39_n109,
         SD1_SB_inst_SD1_SB_bit_inst_39_n108,
         SD1_SB_inst_SD1_SB_bit_inst_39_n107,
         SD1_SB_inst_SD1_SB_bit_inst_39_n106,
         SD1_SB_inst_SD1_SB_bit_inst_39_n105,
         SD1_SB_inst_SD1_SB_bit_inst_39_n104,
         SD1_SB_inst_SD1_SB_bit_inst_39_n103,
         SD1_SB_inst_SD1_SB_bit_inst_39_n102,
         SD1_SB_inst_SD1_SB_bit_inst_39_n101,
         SD1_SB_inst_SD1_SB_bit_inst_39_n100,
         SD1_SB_inst_SD1_SB_bit_inst_40_n131,
         SD1_SB_inst_SD1_SB_bit_inst_40_n130,
         SD1_SB_inst_SD1_SB_bit_inst_40_n129,
         SD1_SB_inst_SD1_SB_bit_inst_40_n128,
         SD1_SB_inst_SD1_SB_bit_inst_40_n127,
         SD1_SB_inst_SD1_SB_bit_inst_40_n126,
         SD1_SB_inst_SD1_SB_bit_inst_40_n125,
         SD1_SB_inst_SD1_SB_bit_inst_40_n124,
         SD1_SB_inst_SD1_SB_bit_inst_40_n123,
         SD1_SB_inst_SD1_SB_bit_inst_40_n122,
         SD1_SB_inst_SD1_SB_bit_inst_40_n121,
         SD1_SB_inst_SD1_SB_bit_inst_40_n120,
         SD1_SB_inst_SD1_SB_bit_inst_40_n119,
         SD1_SB_inst_SD1_SB_bit_inst_40_n118,
         SD1_SB_inst_SD1_SB_bit_inst_40_n117,
         SD1_SB_inst_SD1_SB_bit_inst_40_n116,
         SD1_SB_inst_SD1_SB_bit_inst_40_n115,
         SD1_SB_inst_SD1_SB_bit_inst_40_n114,
         SD1_SB_inst_SD1_SB_bit_inst_40_n113,
         SD1_SB_inst_SD1_SB_bit_inst_40_n112,
         SD1_SB_inst_SD1_SB_bit_inst_40_n111,
         SD1_SB_inst_SD1_SB_bit_inst_40_n110,
         SD1_SB_inst_SD1_SB_bit_inst_40_n109,
         SD1_SB_inst_SD1_SB_bit_inst_40_n108,
         SD1_SB_inst_SD1_SB_bit_inst_40_n107,
         SD1_SB_inst_SD1_SB_bit_inst_40_n106,
         SD1_SB_inst_SD1_SB_bit_inst_40_n105,
         SD1_SB_inst_SD1_SB_bit_inst_40_n104,
         SD1_SB_inst_SD1_SB_bit_inst_40_n103,
         SD1_SB_inst_SD1_SB_bit_inst_40_n102,
         SD1_SB_inst_SD1_SB_bit_inst_40_n101,
         SD1_SB_inst_SD1_SB_bit_inst_40_n100,
         SD1_SB_inst_SD1_SB_bit_inst_40_n99,
         SD1_SB_inst_SD1_SB_bit_inst_40_n98,
         SD1_SB_inst_SD1_SB_bit_inst_40_n97,
         SD1_SB_inst_SD1_SB_bit_inst_40_n96,
         SD1_SB_inst_SD1_SB_bit_inst_40_n95,
         SD1_SB_inst_SD1_SB_bit_inst_40_n94,
         SD1_SB_inst_SD1_SB_bit_inst_40_n93,
         SD1_SB_inst_SD1_SB_bit_inst_40_n92,
         SD1_SB_inst_SD1_SB_bit_inst_41_n110,
         SD1_SB_inst_SD1_SB_bit_inst_41_n109,
         SD1_SB_inst_SD1_SB_bit_inst_41_n108,
         SD1_SB_inst_SD1_SB_bit_inst_41_n107,
         SD1_SB_inst_SD1_SB_bit_inst_41_n106,
         SD1_SB_inst_SD1_SB_bit_inst_41_n105,
         SD1_SB_inst_SD1_SB_bit_inst_41_n104,
         SD1_SB_inst_SD1_SB_bit_inst_41_n103,
         SD1_SB_inst_SD1_SB_bit_inst_41_n102,
         SD1_SB_inst_SD1_SB_bit_inst_41_n101,
         SD1_SB_inst_SD1_SB_bit_inst_41_n100,
         SD1_SB_inst_SD1_SB_bit_inst_41_n99,
         SD1_SB_inst_SD1_SB_bit_inst_41_n98,
         SD1_SB_inst_SD1_SB_bit_inst_41_n97,
         SD1_SB_inst_SD1_SB_bit_inst_41_n96,
         SD1_SB_inst_SD1_SB_bit_inst_41_n95,
         SD1_SB_inst_SD1_SB_bit_inst_41_n94,
         SD1_SB_inst_SD1_SB_bit_inst_41_n93,
         SD1_SB_inst_SD1_SB_bit_inst_41_n92,
         SD1_SB_inst_SD1_SB_bit_inst_41_n91,
         SD1_SB_inst_SD1_SB_bit_inst_41_n90,
         SD1_SB_inst_SD1_SB_bit_inst_41_n89,
         SD1_SB_inst_SD1_SB_bit_inst_41_n88,
         SD1_SB_inst_SD1_SB_bit_inst_41_n87,
         SD1_SB_inst_SD1_SB_bit_inst_41_n86,
         SD1_SB_inst_SD1_SB_bit_inst_41_n85,
         SD1_SB_inst_SD1_SB_bit_inst_41_n84,
         SD1_SB_inst_SD1_SB_bit_inst_41_n83,
         SD1_SB_inst_SD1_SB_bit_inst_41_n82,
         SD1_SB_inst_SD1_SB_bit_inst_41_n81,
         SD1_SB_inst_SD1_SB_bit_inst_41_n80,
         SD1_SB_inst_SD1_SB_bit_inst_41_n79,
         SD1_SB_inst_SD1_SB_bit_inst_41_n78,
         SD1_SB_inst_SD1_SB_bit_inst_41_n77,
         SD1_SB_inst_SD1_SB_bit_inst_42_n138,
         SD1_SB_inst_SD1_SB_bit_inst_42_n137,
         SD1_SB_inst_SD1_SB_bit_inst_42_n136,
         SD1_SB_inst_SD1_SB_bit_inst_42_n135,
         SD1_SB_inst_SD1_SB_bit_inst_42_n134,
         SD1_SB_inst_SD1_SB_bit_inst_42_n133,
         SD1_SB_inst_SD1_SB_bit_inst_42_n132,
         SD1_SB_inst_SD1_SB_bit_inst_42_n131,
         SD1_SB_inst_SD1_SB_bit_inst_42_n130,
         SD1_SB_inst_SD1_SB_bit_inst_42_n129,
         SD1_SB_inst_SD1_SB_bit_inst_42_n128,
         SD1_SB_inst_SD1_SB_bit_inst_42_n127,
         SD1_SB_inst_SD1_SB_bit_inst_42_n126,
         SD1_SB_inst_SD1_SB_bit_inst_42_n125,
         SD1_SB_inst_SD1_SB_bit_inst_42_n124,
         SD1_SB_inst_SD1_SB_bit_inst_42_n123,
         SD1_SB_inst_SD1_SB_bit_inst_42_n122,
         SD1_SB_inst_SD1_SB_bit_inst_42_n121,
         SD1_SB_inst_SD1_SB_bit_inst_42_n120,
         SD1_SB_inst_SD1_SB_bit_inst_42_n119,
         SD1_SB_inst_SD1_SB_bit_inst_42_n118,
         SD1_SB_inst_SD1_SB_bit_inst_42_n117,
         SD1_SB_inst_SD1_SB_bit_inst_42_n116,
         SD1_SB_inst_SD1_SB_bit_inst_42_n115,
         SD1_SB_inst_SD1_SB_bit_inst_42_n114,
         SD1_SB_inst_SD1_SB_bit_inst_42_n113,
         SD1_SB_inst_SD1_SB_bit_inst_42_n112,
         SD1_SB_inst_SD1_SB_bit_inst_42_n111,
         SD1_SB_inst_SD1_SB_bit_inst_42_n110,
         SD1_SB_inst_SD1_SB_bit_inst_42_n109,
         SD1_SB_inst_SD1_SB_bit_inst_42_n108,
         SD1_SB_inst_SD1_SB_bit_inst_42_n107,
         SD1_SB_inst_SD1_SB_bit_inst_42_n106,
         SD1_SB_inst_SD1_SB_bit_inst_42_n105,
         SD1_SB_inst_SD1_SB_bit_inst_42_n104,
         SD1_SB_inst_SD1_SB_bit_inst_42_n103,
         SD1_SB_inst_SD1_SB_bit_inst_42_n102,
         SD1_SB_inst_SD1_SB_bit_inst_42_n101,
         SD1_SB_inst_SD1_SB_bit_inst_42_n100,
         SD1_SB_inst_SD1_SB_bit_inst_42_n99,
         SD1_SB_inst_SD1_SB_bit_inst_42_n98,
         SD1_SB_inst_SD1_SB_bit_inst_42_n97,
         SD1_SB_inst_SD1_SB_bit_inst_43_n141,
         SD1_SB_inst_SD1_SB_bit_inst_43_n140,
         SD1_SB_inst_SD1_SB_bit_inst_43_n139,
         SD1_SB_inst_SD1_SB_bit_inst_43_n138,
         SD1_SB_inst_SD1_SB_bit_inst_43_n137,
         SD1_SB_inst_SD1_SB_bit_inst_43_n136,
         SD1_SB_inst_SD1_SB_bit_inst_43_n135,
         SD1_SB_inst_SD1_SB_bit_inst_43_n134,
         SD1_SB_inst_SD1_SB_bit_inst_43_n133,
         SD1_SB_inst_SD1_SB_bit_inst_43_n132,
         SD1_SB_inst_SD1_SB_bit_inst_43_n131,
         SD1_SB_inst_SD1_SB_bit_inst_43_n130,
         SD1_SB_inst_SD1_SB_bit_inst_43_n129,
         SD1_SB_inst_SD1_SB_bit_inst_43_n128,
         SD1_SB_inst_SD1_SB_bit_inst_43_n127,
         SD1_SB_inst_SD1_SB_bit_inst_43_n126,
         SD1_SB_inst_SD1_SB_bit_inst_43_n125,
         SD1_SB_inst_SD1_SB_bit_inst_43_n124,
         SD1_SB_inst_SD1_SB_bit_inst_43_n123,
         SD1_SB_inst_SD1_SB_bit_inst_43_n122,
         SD1_SB_inst_SD1_SB_bit_inst_43_n121,
         SD1_SB_inst_SD1_SB_bit_inst_43_n120,
         SD1_SB_inst_SD1_SB_bit_inst_43_n119,
         SD1_SB_inst_SD1_SB_bit_inst_43_n118,
         SD1_SB_inst_SD1_SB_bit_inst_43_n117,
         SD1_SB_inst_SD1_SB_bit_inst_43_n116,
         SD1_SB_inst_SD1_SB_bit_inst_43_n115,
         SD1_SB_inst_SD1_SB_bit_inst_43_n114,
         SD1_SB_inst_SD1_SB_bit_inst_43_n113,
         SD1_SB_inst_SD1_SB_bit_inst_43_n112,
         SD1_SB_inst_SD1_SB_bit_inst_43_n111,
         SD1_SB_inst_SD1_SB_bit_inst_43_n110,
         SD1_SB_inst_SD1_SB_bit_inst_43_n109,
         SD1_SB_inst_SD1_SB_bit_inst_43_n108,
         SD1_SB_inst_SD1_SB_bit_inst_43_n107,
         SD1_SB_inst_SD1_SB_bit_inst_43_n106,
         SD1_SB_inst_SD1_SB_bit_inst_43_n105,
         SD1_SB_inst_SD1_SB_bit_inst_43_n104,
         SD1_SB_inst_SD1_SB_bit_inst_43_n103,
         SD1_SB_inst_SD1_SB_bit_inst_43_n102,
         SD1_SB_inst_SD1_SB_bit_inst_43_n101,
         SD1_SB_inst_SD1_SB_bit_inst_43_n100,
         SD1_SB_inst_SD1_SB_bit_inst_44_n131,
         SD1_SB_inst_SD1_SB_bit_inst_44_n130,
         SD1_SB_inst_SD1_SB_bit_inst_44_n129,
         SD1_SB_inst_SD1_SB_bit_inst_44_n128,
         SD1_SB_inst_SD1_SB_bit_inst_44_n127,
         SD1_SB_inst_SD1_SB_bit_inst_44_n126,
         SD1_SB_inst_SD1_SB_bit_inst_44_n125,
         SD1_SB_inst_SD1_SB_bit_inst_44_n124,
         SD1_SB_inst_SD1_SB_bit_inst_44_n123,
         SD1_SB_inst_SD1_SB_bit_inst_44_n122,
         SD1_SB_inst_SD1_SB_bit_inst_44_n121,
         SD1_SB_inst_SD1_SB_bit_inst_44_n120,
         SD1_SB_inst_SD1_SB_bit_inst_44_n119,
         SD1_SB_inst_SD1_SB_bit_inst_44_n118,
         SD1_SB_inst_SD1_SB_bit_inst_44_n117,
         SD1_SB_inst_SD1_SB_bit_inst_44_n116,
         SD1_SB_inst_SD1_SB_bit_inst_44_n115,
         SD1_SB_inst_SD1_SB_bit_inst_44_n114,
         SD1_SB_inst_SD1_SB_bit_inst_44_n113,
         SD1_SB_inst_SD1_SB_bit_inst_44_n112,
         SD1_SB_inst_SD1_SB_bit_inst_44_n111,
         SD1_SB_inst_SD1_SB_bit_inst_44_n110,
         SD1_SB_inst_SD1_SB_bit_inst_44_n109,
         SD1_SB_inst_SD1_SB_bit_inst_44_n108,
         SD1_SB_inst_SD1_SB_bit_inst_44_n107,
         SD1_SB_inst_SD1_SB_bit_inst_44_n106,
         SD1_SB_inst_SD1_SB_bit_inst_44_n105,
         SD1_SB_inst_SD1_SB_bit_inst_44_n104,
         SD1_SB_inst_SD1_SB_bit_inst_44_n103,
         SD1_SB_inst_SD1_SB_bit_inst_44_n102,
         SD1_SB_inst_SD1_SB_bit_inst_44_n101,
         SD1_SB_inst_SD1_SB_bit_inst_44_n100,
         SD1_SB_inst_SD1_SB_bit_inst_44_n99,
         SD1_SB_inst_SD1_SB_bit_inst_44_n98,
         SD1_SB_inst_SD1_SB_bit_inst_44_n97,
         SD1_SB_inst_SD1_SB_bit_inst_44_n96,
         SD1_SB_inst_SD1_SB_bit_inst_44_n95,
         SD1_SB_inst_SD1_SB_bit_inst_44_n94,
         SD1_SB_inst_SD1_SB_bit_inst_44_n93,
         SD1_SB_inst_SD1_SB_bit_inst_44_n92,
         SD1_SB_inst_SD1_SB_bit_inst_45_n110,
         SD1_SB_inst_SD1_SB_bit_inst_45_n109,
         SD1_SB_inst_SD1_SB_bit_inst_45_n108,
         SD1_SB_inst_SD1_SB_bit_inst_45_n107,
         SD1_SB_inst_SD1_SB_bit_inst_45_n106,
         SD1_SB_inst_SD1_SB_bit_inst_45_n105,
         SD1_SB_inst_SD1_SB_bit_inst_45_n104,
         SD1_SB_inst_SD1_SB_bit_inst_45_n103,
         SD1_SB_inst_SD1_SB_bit_inst_45_n102,
         SD1_SB_inst_SD1_SB_bit_inst_45_n101,
         SD1_SB_inst_SD1_SB_bit_inst_45_n100,
         SD1_SB_inst_SD1_SB_bit_inst_45_n99,
         SD1_SB_inst_SD1_SB_bit_inst_45_n98,
         SD1_SB_inst_SD1_SB_bit_inst_45_n97,
         SD1_SB_inst_SD1_SB_bit_inst_45_n96,
         SD1_SB_inst_SD1_SB_bit_inst_45_n95,
         SD1_SB_inst_SD1_SB_bit_inst_45_n94,
         SD1_SB_inst_SD1_SB_bit_inst_45_n93,
         SD1_SB_inst_SD1_SB_bit_inst_45_n92,
         SD1_SB_inst_SD1_SB_bit_inst_45_n91,
         SD1_SB_inst_SD1_SB_bit_inst_45_n90,
         SD1_SB_inst_SD1_SB_bit_inst_45_n89,
         SD1_SB_inst_SD1_SB_bit_inst_45_n88,
         SD1_SB_inst_SD1_SB_bit_inst_45_n87,
         SD1_SB_inst_SD1_SB_bit_inst_45_n86,
         SD1_SB_inst_SD1_SB_bit_inst_45_n85,
         SD1_SB_inst_SD1_SB_bit_inst_45_n84,
         SD1_SB_inst_SD1_SB_bit_inst_45_n83,
         SD1_SB_inst_SD1_SB_bit_inst_45_n82,
         SD1_SB_inst_SD1_SB_bit_inst_45_n81,
         SD1_SB_inst_SD1_SB_bit_inst_45_n80,
         SD1_SB_inst_SD1_SB_bit_inst_45_n79,
         SD1_SB_inst_SD1_SB_bit_inst_45_n78,
         SD1_SB_inst_SD1_SB_bit_inst_45_n77,
         SD1_SB_inst_SD1_SB_bit_inst_46_n138,
         SD1_SB_inst_SD1_SB_bit_inst_46_n137,
         SD1_SB_inst_SD1_SB_bit_inst_46_n136,
         SD1_SB_inst_SD1_SB_bit_inst_46_n135,
         SD1_SB_inst_SD1_SB_bit_inst_46_n134,
         SD1_SB_inst_SD1_SB_bit_inst_46_n133,
         SD1_SB_inst_SD1_SB_bit_inst_46_n132,
         SD1_SB_inst_SD1_SB_bit_inst_46_n131,
         SD1_SB_inst_SD1_SB_bit_inst_46_n130,
         SD1_SB_inst_SD1_SB_bit_inst_46_n129,
         SD1_SB_inst_SD1_SB_bit_inst_46_n128,
         SD1_SB_inst_SD1_SB_bit_inst_46_n127,
         SD1_SB_inst_SD1_SB_bit_inst_46_n126,
         SD1_SB_inst_SD1_SB_bit_inst_46_n125,
         SD1_SB_inst_SD1_SB_bit_inst_46_n124,
         SD1_SB_inst_SD1_SB_bit_inst_46_n123,
         SD1_SB_inst_SD1_SB_bit_inst_46_n122,
         SD1_SB_inst_SD1_SB_bit_inst_46_n121,
         SD1_SB_inst_SD1_SB_bit_inst_46_n120,
         SD1_SB_inst_SD1_SB_bit_inst_46_n119,
         SD1_SB_inst_SD1_SB_bit_inst_46_n118,
         SD1_SB_inst_SD1_SB_bit_inst_46_n117,
         SD1_SB_inst_SD1_SB_bit_inst_46_n116,
         SD1_SB_inst_SD1_SB_bit_inst_46_n115,
         SD1_SB_inst_SD1_SB_bit_inst_46_n114,
         SD1_SB_inst_SD1_SB_bit_inst_46_n113,
         SD1_SB_inst_SD1_SB_bit_inst_46_n112,
         SD1_SB_inst_SD1_SB_bit_inst_46_n111,
         SD1_SB_inst_SD1_SB_bit_inst_46_n110,
         SD1_SB_inst_SD1_SB_bit_inst_46_n109,
         SD1_SB_inst_SD1_SB_bit_inst_46_n108,
         SD1_SB_inst_SD1_SB_bit_inst_46_n107,
         SD1_SB_inst_SD1_SB_bit_inst_46_n106,
         SD1_SB_inst_SD1_SB_bit_inst_46_n105,
         SD1_SB_inst_SD1_SB_bit_inst_46_n104,
         SD1_SB_inst_SD1_SB_bit_inst_46_n103,
         SD1_SB_inst_SD1_SB_bit_inst_46_n102,
         SD1_SB_inst_SD1_SB_bit_inst_46_n101,
         SD1_SB_inst_SD1_SB_bit_inst_46_n100,
         SD1_SB_inst_SD1_SB_bit_inst_46_n99,
         SD1_SB_inst_SD1_SB_bit_inst_46_n98,
         SD1_SB_inst_SD1_SB_bit_inst_46_n97,
         SD1_SB_inst_SD1_SB_bit_inst_47_n141,
         SD1_SB_inst_SD1_SB_bit_inst_47_n140,
         SD1_SB_inst_SD1_SB_bit_inst_47_n139,
         SD1_SB_inst_SD1_SB_bit_inst_47_n138,
         SD1_SB_inst_SD1_SB_bit_inst_47_n137,
         SD1_SB_inst_SD1_SB_bit_inst_47_n136,
         SD1_SB_inst_SD1_SB_bit_inst_47_n135,
         SD1_SB_inst_SD1_SB_bit_inst_47_n134,
         SD1_SB_inst_SD1_SB_bit_inst_47_n133,
         SD1_SB_inst_SD1_SB_bit_inst_47_n132,
         SD1_SB_inst_SD1_SB_bit_inst_47_n131,
         SD1_SB_inst_SD1_SB_bit_inst_47_n130,
         SD1_SB_inst_SD1_SB_bit_inst_47_n129,
         SD1_SB_inst_SD1_SB_bit_inst_47_n128,
         SD1_SB_inst_SD1_SB_bit_inst_47_n127,
         SD1_SB_inst_SD1_SB_bit_inst_47_n126,
         SD1_SB_inst_SD1_SB_bit_inst_47_n125,
         SD1_SB_inst_SD1_SB_bit_inst_47_n124,
         SD1_SB_inst_SD1_SB_bit_inst_47_n123,
         SD1_SB_inst_SD1_SB_bit_inst_47_n122,
         SD1_SB_inst_SD1_SB_bit_inst_47_n121,
         SD1_SB_inst_SD1_SB_bit_inst_47_n120,
         SD1_SB_inst_SD1_SB_bit_inst_47_n119,
         SD1_SB_inst_SD1_SB_bit_inst_47_n118,
         SD1_SB_inst_SD1_SB_bit_inst_47_n117,
         SD1_SB_inst_SD1_SB_bit_inst_47_n116,
         SD1_SB_inst_SD1_SB_bit_inst_47_n115,
         SD1_SB_inst_SD1_SB_bit_inst_47_n114,
         SD1_SB_inst_SD1_SB_bit_inst_47_n113,
         SD1_SB_inst_SD1_SB_bit_inst_47_n112,
         SD1_SB_inst_SD1_SB_bit_inst_47_n111,
         SD1_SB_inst_SD1_SB_bit_inst_47_n110,
         SD1_SB_inst_SD1_SB_bit_inst_47_n109,
         SD1_SB_inst_SD1_SB_bit_inst_47_n108,
         SD1_SB_inst_SD1_SB_bit_inst_47_n107,
         SD1_SB_inst_SD1_SB_bit_inst_47_n106,
         SD1_SB_inst_SD1_SB_bit_inst_47_n105,
         SD1_SB_inst_SD1_SB_bit_inst_47_n104,
         SD1_SB_inst_SD1_SB_bit_inst_47_n103,
         SD1_SB_inst_SD1_SB_bit_inst_47_n102,
         SD1_SB_inst_SD1_SB_bit_inst_47_n101,
         SD1_SB_inst_SD1_SB_bit_inst_47_n100,
         SD1_SB_inst_SD1_SB_bit_inst_48_n131,
         SD1_SB_inst_SD1_SB_bit_inst_48_n130,
         SD1_SB_inst_SD1_SB_bit_inst_48_n129,
         SD1_SB_inst_SD1_SB_bit_inst_48_n128,
         SD1_SB_inst_SD1_SB_bit_inst_48_n127,
         SD1_SB_inst_SD1_SB_bit_inst_48_n126,
         SD1_SB_inst_SD1_SB_bit_inst_48_n125,
         SD1_SB_inst_SD1_SB_bit_inst_48_n124,
         SD1_SB_inst_SD1_SB_bit_inst_48_n123,
         SD1_SB_inst_SD1_SB_bit_inst_48_n122,
         SD1_SB_inst_SD1_SB_bit_inst_48_n121,
         SD1_SB_inst_SD1_SB_bit_inst_48_n120,
         SD1_SB_inst_SD1_SB_bit_inst_48_n119,
         SD1_SB_inst_SD1_SB_bit_inst_48_n118,
         SD1_SB_inst_SD1_SB_bit_inst_48_n117,
         SD1_SB_inst_SD1_SB_bit_inst_48_n116,
         SD1_SB_inst_SD1_SB_bit_inst_48_n115,
         SD1_SB_inst_SD1_SB_bit_inst_48_n114,
         SD1_SB_inst_SD1_SB_bit_inst_48_n113,
         SD1_SB_inst_SD1_SB_bit_inst_48_n112,
         SD1_SB_inst_SD1_SB_bit_inst_48_n111,
         SD1_SB_inst_SD1_SB_bit_inst_48_n110,
         SD1_SB_inst_SD1_SB_bit_inst_48_n109,
         SD1_SB_inst_SD1_SB_bit_inst_48_n108,
         SD1_SB_inst_SD1_SB_bit_inst_48_n107,
         SD1_SB_inst_SD1_SB_bit_inst_48_n106,
         SD1_SB_inst_SD1_SB_bit_inst_48_n105,
         SD1_SB_inst_SD1_SB_bit_inst_48_n104,
         SD1_SB_inst_SD1_SB_bit_inst_48_n103,
         SD1_SB_inst_SD1_SB_bit_inst_48_n102,
         SD1_SB_inst_SD1_SB_bit_inst_48_n101,
         SD1_SB_inst_SD1_SB_bit_inst_48_n100,
         SD1_SB_inst_SD1_SB_bit_inst_48_n99,
         SD1_SB_inst_SD1_SB_bit_inst_48_n98,
         SD1_SB_inst_SD1_SB_bit_inst_48_n97,
         SD1_SB_inst_SD1_SB_bit_inst_48_n96,
         SD1_SB_inst_SD1_SB_bit_inst_48_n95,
         SD1_SB_inst_SD1_SB_bit_inst_48_n94,
         SD1_SB_inst_SD1_SB_bit_inst_48_n93,
         SD1_SB_inst_SD1_SB_bit_inst_48_n92,
         SD1_SB_inst_SD1_SB_bit_inst_49_n110,
         SD1_SB_inst_SD1_SB_bit_inst_49_n109,
         SD1_SB_inst_SD1_SB_bit_inst_49_n108,
         SD1_SB_inst_SD1_SB_bit_inst_49_n107,
         SD1_SB_inst_SD1_SB_bit_inst_49_n106,
         SD1_SB_inst_SD1_SB_bit_inst_49_n105,
         SD1_SB_inst_SD1_SB_bit_inst_49_n104,
         SD1_SB_inst_SD1_SB_bit_inst_49_n103,
         SD1_SB_inst_SD1_SB_bit_inst_49_n102,
         SD1_SB_inst_SD1_SB_bit_inst_49_n101,
         SD1_SB_inst_SD1_SB_bit_inst_49_n100,
         SD1_SB_inst_SD1_SB_bit_inst_49_n99,
         SD1_SB_inst_SD1_SB_bit_inst_49_n98,
         SD1_SB_inst_SD1_SB_bit_inst_49_n97,
         SD1_SB_inst_SD1_SB_bit_inst_49_n96,
         SD1_SB_inst_SD1_SB_bit_inst_49_n95,
         SD1_SB_inst_SD1_SB_bit_inst_49_n94,
         SD1_SB_inst_SD1_SB_bit_inst_49_n93,
         SD1_SB_inst_SD1_SB_bit_inst_49_n92,
         SD1_SB_inst_SD1_SB_bit_inst_49_n91,
         SD1_SB_inst_SD1_SB_bit_inst_49_n90,
         SD1_SB_inst_SD1_SB_bit_inst_49_n89,
         SD1_SB_inst_SD1_SB_bit_inst_49_n88,
         SD1_SB_inst_SD1_SB_bit_inst_49_n87,
         SD1_SB_inst_SD1_SB_bit_inst_49_n86,
         SD1_SB_inst_SD1_SB_bit_inst_49_n85,
         SD1_SB_inst_SD1_SB_bit_inst_49_n84,
         SD1_SB_inst_SD1_SB_bit_inst_49_n83,
         SD1_SB_inst_SD1_SB_bit_inst_49_n82,
         SD1_SB_inst_SD1_SB_bit_inst_49_n81,
         SD1_SB_inst_SD1_SB_bit_inst_49_n80,
         SD1_SB_inst_SD1_SB_bit_inst_49_n79,
         SD1_SB_inst_SD1_SB_bit_inst_49_n78,
         SD1_SB_inst_SD1_SB_bit_inst_49_n77,
         SD1_SB_inst_SD1_SB_bit_inst_50_n138,
         SD1_SB_inst_SD1_SB_bit_inst_50_n137,
         SD1_SB_inst_SD1_SB_bit_inst_50_n136,
         SD1_SB_inst_SD1_SB_bit_inst_50_n135,
         SD1_SB_inst_SD1_SB_bit_inst_50_n134,
         SD1_SB_inst_SD1_SB_bit_inst_50_n133,
         SD1_SB_inst_SD1_SB_bit_inst_50_n132,
         SD1_SB_inst_SD1_SB_bit_inst_50_n131,
         SD1_SB_inst_SD1_SB_bit_inst_50_n130,
         SD1_SB_inst_SD1_SB_bit_inst_50_n129,
         SD1_SB_inst_SD1_SB_bit_inst_50_n128,
         SD1_SB_inst_SD1_SB_bit_inst_50_n127,
         SD1_SB_inst_SD1_SB_bit_inst_50_n126,
         SD1_SB_inst_SD1_SB_bit_inst_50_n125,
         SD1_SB_inst_SD1_SB_bit_inst_50_n124,
         SD1_SB_inst_SD1_SB_bit_inst_50_n123,
         SD1_SB_inst_SD1_SB_bit_inst_50_n122,
         SD1_SB_inst_SD1_SB_bit_inst_50_n121,
         SD1_SB_inst_SD1_SB_bit_inst_50_n120,
         SD1_SB_inst_SD1_SB_bit_inst_50_n119,
         SD1_SB_inst_SD1_SB_bit_inst_50_n118,
         SD1_SB_inst_SD1_SB_bit_inst_50_n117,
         SD1_SB_inst_SD1_SB_bit_inst_50_n116,
         SD1_SB_inst_SD1_SB_bit_inst_50_n115,
         SD1_SB_inst_SD1_SB_bit_inst_50_n114,
         SD1_SB_inst_SD1_SB_bit_inst_50_n113,
         SD1_SB_inst_SD1_SB_bit_inst_50_n112,
         SD1_SB_inst_SD1_SB_bit_inst_50_n111,
         SD1_SB_inst_SD1_SB_bit_inst_50_n110,
         SD1_SB_inst_SD1_SB_bit_inst_50_n109,
         SD1_SB_inst_SD1_SB_bit_inst_50_n108,
         SD1_SB_inst_SD1_SB_bit_inst_50_n107,
         SD1_SB_inst_SD1_SB_bit_inst_50_n106,
         SD1_SB_inst_SD1_SB_bit_inst_50_n105,
         SD1_SB_inst_SD1_SB_bit_inst_50_n104,
         SD1_SB_inst_SD1_SB_bit_inst_50_n103,
         SD1_SB_inst_SD1_SB_bit_inst_50_n102,
         SD1_SB_inst_SD1_SB_bit_inst_50_n101,
         SD1_SB_inst_SD1_SB_bit_inst_50_n100,
         SD1_SB_inst_SD1_SB_bit_inst_50_n99,
         SD1_SB_inst_SD1_SB_bit_inst_50_n98,
         SD1_SB_inst_SD1_SB_bit_inst_50_n97,
         SD1_SB_inst_SD1_SB_bit_inst_51_n141,
         SD1_SB_inst_SD1_SB_bit_inst_51_n140,
         SD1_SB_inst_SD1_SB_bit_inst_51_n139,
         SD1_SB_inst_SD1_SB_bit_inst_51_n138,
         SD1_SB_inst_SD1_SB_bit_inst_51_n137,
         SD1_SB_inst_SD1_SB_bit_inst_51_n136,
         SD1_SB_inst_SD1_SB_bit_inst_51_n135,
         SD1_SB_inst_SD1_SB_bit_inst_51_n134,
         SD1_SB_inst_SD1_SB_bit_inst_51_n133,
         SD1_SB_inst_SD1_SB_bit_inst_51_n132,
         SD1_SB_inst_SD1_SB_bit_inst_51_n131,
         SD1_SB_inst_SD1_SB_bit_inst_51_n130,
         SD1_SB_inst_SD1_SB_bit_inst_51_n129,
         SD1_SB_inst_SD1_SB_bit_inst_51_n128,
         SD1_SB_inst_SD1_SB_bit_inst_51_n127,
         SD1_SB_inst_SD1_SB_bit_inst_51_n126,
         SD1_SB_inst_SD1_SB_bit_inst_51_n125,
         SD1_SB_inst_SD1_SB_bit_inst_51_n124,
         SD1_SB_inst_SD1_SB_bit_inst_51_n123,
         SD1_SB_inst_SD1_SB_bit_inst_51_n122,
         SD1_SB_inst_SD1_SB_bit_inst_51_n121,
         SD1_SB_inst_SD1_SB_bit_inst_51_n120,
         SD1_SB_inst_SD1_SB_bit_inst_51_n119,
         SD1_SB_inst_SD1_SB_bit_inst_51_n118,
         SD1_SB_inst_SD1_SB_bit_inst_51_n117,
         SD1_SB_inst_SD1_SB_bit_inst_51_n116,
         SD1_SB_inst_SD1_SB_bit_inst_51_n115,
         SD1_SB_inst_SD1_SB_bit_inst_51_n114,
         SD1_SB_inst_SD1_SB_bit_inst_51_n113,
         SD1_SB_inst_SD1_SB_bit_inst_51_n112,
         SD1_SB_inst_SD1_SB_bit_inst_51_n111,
         SD1_SB_inst_SD1_SB_bit_inst_51_n110,
         SD1_SB_inst_SD1_SB_bit_inst_51_n109,
         SD1_SB_inst_SD1_SB_bit_inst_51_n108,
         SD1_SB_inst_SD1_SB_bit_inst_51_n107,
         SD1_SB_inst_SD1_SB_bit_inst_51_n106,
         SD1_SB_inst_SD1_SB_bit_inst_51_n105,
         SD1_SB_inst_SD1_SB_bit_inst_51_n104,
         SD1_SB_inst_SD1_SB_bit_inst_51_n103,
         SD1_SB_inst_SD1_SB_bit_inst_51_n102,
         SD1_SB_inst_SD1_SB_bit_inst_51_n101,
         SD1_SB_inst_SD1_SB_bit_inst_51_n100,
         SD1_SB_inst_SD1_SB_bit_inst_52_n131,
         SD1_SB_inst_SD1_SB_bit_inst_52_n130,
         SD1_SB_inst_SD1_SB_bit_inst_52_n129,
         SD1_SB_inst_SD1_SB_bit_inst_52_n128,
         SD1_SB_inst_SD1_SB_bit_inst_52_n127,
         SD1_SB_inst_SD1_SB_bit_inst_52_n126,
         SD1_SB_inst_SD1_SB_bit_inst_52_n125,
         SD1_SB_inst_SD1_SB_bit_inst_52_n124,
         SD1_SB_inst_SD1_SB_bit_inst_52_n123,
         SD1_SB_inst_SD1_SB_bit_inst_52_n122,
         SD1_SB_inst_SD1_SB_bit_inst_52_n121,
         SD1_SB_inst_SD1_SB_bit_inst_52_n120,
         SD1_SB_inst_SD1_SB_bit_inst_52_n119,
         SD1_SB_inst_SD1_SB_bit_inst_52_n118,
         SD1_SB_inst_SD1_SB_bit_inst_52_n117,
         SD1_SB_inst_SD1_SB_bit_inst_52_n116,
         SD1_SB_inst_SD1_SB_bit_inst_52_n115,
         SD1_SB_inst_SD1_SB_bit_inst_52_n114,
         SD1_SB_inst_SD1_SB_bit_inst_52_n113,
         SD1_SB_inst_SD1_SB_bit_inst_52_n112,
         SD1_SB_inst_SD1_SB_bit_inst_52_n111,
         SD1_SB_inst_SD1_SB_bit_inst_52_n110,
         SD1_SB_inst_SD1_SB_bit_inst_52_n109,
         SD1_SB_inst_SD1_SB_bit_inst_52_n108,
         SD1_SB_inst_SD1_SB_bit_inst_52_n107,
         SD1_SB_inst_SD1_SB_bit_inst_52_n106,
         SD1_SB_inst_SD1_SB_bit_inst_52_n105,
         SD1_SB_inst_SD1_SB_bit_inst_52_n104,
         SD1_SB_inst_SD1_SB_bit_inst_52_n103,
         SD1_SB_inst_SD1_SB_bit_inst_52_n102,
         SD1_SB_inst_SD1_SB_bit_inst_52_n101,
         SD1_SB_inst_SD1_SB_bit_inst_52_n100,
         SD1_SB_inst_SD1_SB_bit_inst_52_n99,
         SD1_SB_inst_SD1_SB_bit_inst_52_n98,
         SD1_SB_inst_SD1_SB_bit_inst_52_n97,
         SD1_SB_inst_SD1_SB_bit_inst_52_n96,
         SD1_SB_inst_SD1_SB_bit_inst_52_n95,
         SD1_SB_inst_SD1_SB_bit_inst_52_n94,
         SD1_SB_inst_SD1_SB_bit_inst_52_n93,
         SD1_SB_inst_SD1_SB_bit_inst_52_n92,
         SD1_SB_inst_SD1_SB_bit_inst_53_n110,
         SD1_SB_inst_SD1_SB_bit_inst_53_n109,
         SD1_SB_inst_SD1_SB_bit_inst_53_n108,
         SD1_SB_inst_SD1_SB_bit_inst_53_n107,
         SD1_SB_inst_SD1_SB_bit_inst_53_n106,
         SD1_SB_inst_SD1_SB_bit_inst_53_n105,
         SD1_SB_inst_SD1_SB_bit_inst_53_n104,
         SD1_SB_inst_SD1_SB_bit_inst_53_n103,
         SD1_SB_inst_SD1_SB_bit_inst_53_n102,
         SD1_SB_inst_SD1_SB_bit_inst_53_n101,
         SD1_SB_inst_SD1_SB_bit_inst_53_n100,
         SD1_SB_inst_SD1_SB_bit_inst_53_n99,
         SD1_SB_inst_SD1_SB_bit_inst_53_n98,
         SD1_SB_inst_SD1_SB_bit_inst_53_n97,
         SD1_SB_inst_SD1_SB_bit_inst_53_n96,
         SD1_SB_inst_SD1_SB_bit_inst_53_n95,
         SD1_SB_inst_SD1_SB_bit_inst_53_n94,
         SD1_SB_inst_SD1_SB_bit_inst_53_n93,
         SD1_SB_inst_SD1_SB_bit_inst_53_n92,
         SD1_SB_inst_SD1_SB_bit_inst_53_n91,
         SD1_SB_inst_SD1_SB_bit_inst_53_n90,
         SD1_SB_inst_SD1_SB_bit_inst_53_n89,
         SD1_SB_inst_SD1_SB_bit_inst_53_n88,
         SD1_SB_inst_SD1_SB_bit_inst_53_n87,
         SD1_SB_inst_SD1_SB_bit_inst_53_n86,
         SD1_SB_inst_SD1_SB_bit_inst_53_n85,
         SD1_SB_inst_SD1_SB_bit_inst_53_n84,
         SD1_SB_inst_SD1_SB_bit_inst_53_n83,
         SD1_SB_inst_SD1_SB_bit_inst_53_n82,
         SD1_SB_inst_SD1_SB_bit_inst_53_n81,
         SD1_SB_inst_SD1_SB_bit_inst_53_n80,
         SD1_SB_inst_SD1_SB_bit_inst_53_n79,
         SD1_SB_inst_SD1_SB_bit_inst_53_n78,
         SD1_SB_inst_SD1_SB_bit_inst_53_n77,
         SD1_SB_inst_SD1_SB_bit_inst_54_n138,
         SD1_SB_inst_SD1_SB_bit_inst_54_n137,
         SD1_SB_inst_SD1_SB_bit_inst_54_n136,
         SD1_SB_inst_SD1_SB_bit_inst_54_n135,
         SD1_SB_inst_SD1_SB_bit_inst_54_n134,
         SD1_SB_inst_SD1_SB_bit_inst_54_n133,
         SD1_SB_inst_SD1_SB_bit_inst_54_n132,
         SD1_SB_inst_SD1_SB_bit_inst_54_n131,
         SD1_SB_inst_SD1_SB_bit_inst_54_n130,
         SD1_SB_inst_SD1_SB_bit_inst_54_n129,
         SD1_SB_inst_SD1_SB_bit_inst_54_n128,
         SD1_SB_inst_SD1_SB_bit_inst_54_n127,
         SD1_SB_inst_SD1_SB_bit_inst_54_n126,
         SD1_SB_inst_SD1_SB_bit_inst_54_n125,
         SD1_SB_inst_SD1_SB_bit_inst_54_n124,
         SD1_SB_inst_SD1_SB_bit_inst_54_n123,
         SD1_SB_inst_SD1_SB_bit_inst_54_n122,
         SD1_SB_inst_SD1_SB_bit_inst_54_n121,
         SD1_SB_inst_SD1_SB_bit_inst_54_n120,
         SD1_SB_inst_SD1_SB_bit_inst_54_n119,
         SD1_SB_inst_SD1_SB_bit_inst_54_n118,
         SD1_SB_inst_SD1_SB_bit_inst_54_n117,
         SD1_SB_inst_SD1_SB_bit_inst_54_n116,
         SD1_SB_inst_SD1_SB_bit_inst_54_n115,
         SD1_SB_inst_SD1_SB_bit_inst_54_n114,
         SD1_SB_inst_SD1_SB_bit_inst_54_n113,
         SD1_SB_inst_SD1_SB_bit_inst_54_n112,
         SD1_SB_inst_SD1_SB_bit_inst_54_n111,
         SD1_SB_inst_SD1_SB_bit_inst_54_n110,
         SD1_SB_inst_SD1_SB_bit_inst_54_n109,
         SD1_SB_inst_SD1_SB_bit_inst_54_n108,
         SD1_SB_inst_SD1_SB_bit_inst_54_n107,
         SD1_SB_inst_SD1_SB_bit_inst_54_n106,
         SD1_SB_inst_SD1_SB_bit_inst_54_n105,
         SD1_SB_inst_SD1_SB_bit_inst_54_n104,
         SD1_SB_inst_SD1_SB_bit_inst_54_n103,
         SD1_SB_inst_SD1_SB_bit_inst_54_n102,
         SD1_SB_inst_SD1_SB_bit_inst_54_n101,
         SD1_SB_inst_SD1_SB_bit_inst_54_n100,
         SD1_SB_inst_SD1_SB_bit_inst_54_n99,
         SD1_SB_inst_SD1_SB_bit_inst_54_n98,
         SD1_SB_inst_SD1_SB_bit_inst_54_n97,
         SD1_SB_inst_SD1_SB_bit_inst_55_n141,
         SD1_SB_inst_SD1_SB_bit_inst_55_n140,
         SD1_SB_inst_SD1_SB_bit_inst_55_n139,
         SD1_SB_inst_SD1_SB_bit_inst_55_n138,
         SD1_SB_inst_SD1_SB_bit_inst_55_n137,
         SD1_SB_inst_SD1_SB_bit_inst_55_n136,
         SD1_SB_inst_SD1_SB_bit_inst_55_n135,
         SD1_SB_inst_SD1_SB_bit_inst_55_n134,
         SD1_SB_inst_SD1_SB_bit_inst_55_n133,
         SD1_SB_inst_SD1_SB_bit_inst_55_n132,
         SD1_SB_inst_SD1_SB_bit_inst_55_n131,
         SD1_SB_inst_SD1_SB_bit_inst_55_n130,
         SD1_SB_inst_SD1_SB_bit_inst_55_n129,
         SD1_SB_inst_SD1_SB_bit_inst_55_n128,
         SD1_SB_inst_SD1_SB_bit_inst_55_n127,
         SD1_SB_inst_SD1_SB_bit_inst_55_n126,
         SD1_SB_inst_SD1_SB_bit_inst_55_n125,
         SD1_SB_inst_SD1_SB_bit_inst_55_n124,
         SD1_SB_inst_SD1_SB_bit_inst_55_n123,
         SD1_SB_inst_SD1_SB_bit_inst_55_n122,
         SD1_SB_inst_SD1_SB_bit_inst_55_n121,
         SD1_SB_inst_SD1_SB_bit_inst_55_n120,
         SD1_SB_inst_SD1_SB_bit_inst_55_n119,
         SD1_SB_inst_SD1_SB_bit_inst_55_n118,
         SD1_SB_inst_SD1_SB_bit_inst_55_n117,
         SD1_SB_inst_SD1_SB_bit_inst_55_n116,
         SD1_SB_inst_SD1_SB_bit_inst_55_n115,
         SD1_SB_inst_SD1_SB_bit_inst_55_n114,
         SD1_SB_inst_SD1_SB_bit_inst_55_n113,
         SD1_SB_inst_SD1_SB_bit_inst_55_n112,
         SD1_SB_inst_SD1_SB_bit_inst_55_n111,
         SD1_SB_inst_SD1_SB_bit_inst_55_n110,
         SD1_SB_inst_SD1_SB_bit_inst_55_n109,
         SD1_SB_inst_SD1_SB_bit_inst_55_n108,
         SD1_SB_inst_SD1_SB_bit_inst_55_n107,
         SD1_SB_inst_SD1_SB_bit_inst_55_n106,
         SD1_SB_inst_SD1_SB_bit_inst_55_n105,
         SD1_SB_inst_SD1_SB_bit_inst_55_n104,
         SD1_SB_inst_SD1_SB_bit_inst_55_n103,
         SD1_SB_inst_SD1_SB_bit_inst_55_n102,
         SD1_SB_inst_SD1_SB_bit_inst_55_n101,
         SD1_SB_inst_SD1_SB_bit_inst_55_n100,
         SD1_SB_inst_SD1_SB_bit_inst_56_n131,
         SD1_SB_inst_SD1_SB_bit_inst_56_n130,
         SD1_SB_inst_SD1_SB_bit_inst_56_n129,
         SD1_SB_inst_SD1_SB_bit_inst_56_n128,
         SD1_SB_inst_SD1_SB_bit_inst_56_n127,
         SD1_SB_inst_SD1_SB_bit_inst_56_n126,
         SD1_SB_inst_SD1_SB_bit_inst_56_n125,
         SD1_SB_inst_SD1_SB_bit_inst_56_n124,
         SD1_SB_inst_SD1_SB_bit_inst_56_n123,
         SD1_SB_inst_SD1_SB_bit_inst_56_n122,
         SD1_SB_inst_SD1_SB_bit_inst_56_n121,
         SD1_SB_inst_SD1_SB_bit_inst_56_n120,
         SD1_SB_inst_SD1_SB_bit_inst_56_n119,
         SD1_SB_inst_SD1_SB_bit_inst_56_n118,
         SD1_SB_inst_SD1_SB_bit_inst_56_n117,
         SD1_SB_inst_SD1_SB_bit_inst_56_n116,
         SD1_SB_inst_SD1_SB_bit_inst_56_n115,
         SD1_SB_inst_SD1_SB_bit_inst_56_n114,
         SD1_SB_inst_SD1_SB_bit_inst_56_n113,
         SD1_SB_inst_SD1_SB_bit_inst_56_n112,
         SD1_SB_inst_SD1_SB_bit_inst_56_n111,
         SD1_SB_inst_SD1_SB_bit_inst_56_n110,
         SD1_SB_inst_SD1_SB_bit_inst_56_n109,
         SD1_SB_inst_SD1_SB_bit_inst_56_n108,
         SD1_SB_inst_SD1_SB_bit_inst_56_n107,
         SD1_SB_inst_SD1_SB_bit_inst_56_n106,
         SD1_SB_inst_SD1_SB_bit_inst_56_n105,
         SD1_SB_inst_SD1_SB_bit_inst_56_n104,
         SD1_SB_inst_SD1_SB_bit_inst_56_n103,
         SD1_SB_inst_SD1_SB_bit_inst_56_n102,
         SD1_SB_inst_SD1_SB_bit_inst_56_n101,
         SD1_SB_inst_SD1_SB_bit_inst_56_n100,
         SD1_SB_inst_SD1_SB_bit_inst_56_n99,
         SD1_SB_inst_SD1_SB_bit_inst_56_n98,
         SD1_SB_inst_SD1_SB_bit_inst_56_n97,
         SD1_SB_inst_SD1_SB_bit_inst_56_n96,
         SD1_SB_inst_SD1_SB_bit_inst_56_n95,
         SD1_SB_inst_SD1_SB_bit_inst_56_n94,
         SD1_SB_inst_SD1_SB_bit_inst_56_n93,
         SD1_SB_inst_SD1_SB_bit_inst_56_n92,
         SD1_SB_inst_SD1_SB_bit_inst_57_n110,
         SD1_SB_inst_SD1_SB_bit_inst_57_n109,
         SD1_SB_inst_SD1_SB_bit_inst_57_n108,
         SD1_SB_inst_SD1_SB_bit_inst_57_n107,
         SD1_SB_inst_SD1_SB_bit_inst_57_n106,
         SD1_SB_inst_SD1_SB_bit_inst_57_n105,
         SD1_SB_inst_SD1_SB_bit_inst_57_n104,
         SD1_SB_inst_SD1_SB_bit_inst_57_n103,
         SD1_SB_inst_SD1_SB_bit_inst_57_n102,
         SD1_SB_inst_SD1_SB_bit_inst_57_n101,
         SD1_SB_inst_SD1_SB_bit_inst_57_n100,
         SD1_SB_inst_SD1_SB_bit_inst_57_n99,
         SD1_SB_inst_SD1_SB_bit_inst_57_n98,
         SD1_SB_inst_SD1_SB_bit_inst_57_n97,
         SD1_SB_inst_SD1_SB_bit_inst_57_n96,
         SD1_SB_inst_SD1_SB_bit_inst_57_n95,
         SD1_SB_inst_SD1_SB_bit_inst_57_n94,
         SD1_SB_inst_SD1_SB_bit_inst_57_n93,
         SD1_SB_inst_SD1_SB_bit_inst_57_n92,
         SD1_SB_inst_SD1_SB_bit_inst_57_n91,
         SD1_SB_inst_SD1_SB_bit_inst_57_n90,
         SD1_SB_inst_SD1_SB_bit_inst_57_n89,
         SD1_SB_inst_SD1_SB_bit_inst_57_n88,
         SD1_SB_inst_SD1_SB_bit_inst_57_n87,
         SD1_SB_inst_SD1_SB_bit_inst_57_n86,
         SD1_SB_inst_SD1_SB_bit_inst_57_n85,
         SD1_SB_inst_SD1_SB_bit_inst_57_n84,
         SD1_SB_inst_SD1_SB_bit_inst_57_n83,
         SD1_SB_inst_SD1_SB_bit_inst_57_n82,
         SD1_SB_inst_SD1_SB_bit_inst_57_n81,
         SD1_SB_inst_SD1_SB_bit_inst_57_n80,
         SD1_SB_inst_SD1_SB_bit_inst_57_n79,
         SD1_SB_inst_SD1_SB_bit_inst_57_n78,
         SD1_SB_inst_SD1_SB_bit_inst_57_n77,
         SD1_SB_inst_SD1_SB_bit_inst_58_n138,
         SD1_SB_inst_SD1_SB_bit_inst_58_n137,
         SD1_SB_inst_SD1_SB_bit_inst_58_n136,
         SD1_SB_inst_SD1_SB_bit_inst_58_n135,
         SD1_SB_inst_SD1_SB_bit_inst_58_n134,
         SD1_SB_inst_SD1_SB_bit_inst_58_n133,
         SD1_SB_inst_SD1_SB_bit_inst_58_n132,
         SD1_SB_inst_SD1_SB_bit_inst_58_n131,
         SD1_SB_inst_SD1_SB_bit_inst_58_n130,
         SD1_SB_inst_SD1_SB_bit_inst_58_n129,
         SD1_SB_inst_SD1_SB_bit_inst_58_n128,
         SD1_SB_inst_SD1_SB_bit_inst_58_n127,
         SD1_SB_inst_SD1_SB_bit_inst_58_n126,
         SD1_SB_inst_SD1_SB_bit_inst_58_n125,
         SD1_SB_inst_SD1_SB_bit_inst_58_n124,
         SD1_SB_inst_SD1_SB_bit_inst_58_n123,
         SD1_SB_inst_SD1_SB_bit_inst_58_n122,
         SD1_SB_inst_SD1_SB_bit_inst_58_n121,
         SD1_SB_inst_SD1_SB_bit_inst_58_n120,
         SD1_SB_inst_SD1_SB_bit_inst_58_n119,
         SD1_SB_inst_SD1_SB_bit_inst_58_n118,
         SD1_SB_inst_SD1_SB_bit_inst_58_n117,
         SD1_SB_inst_SD1_SB_bit_inst_58_n116,
         SD1_SB_inst_SD1_SB_bit_inst_58_n115,
         SD1_SB_inst_SD1_SB_bit_inst_58_n114,
         SD1_SB_inst_SD1_SB_bit_inst_58_n113,
         SD1_SB_inst_SD1_SB_bit_inst_58_n112,
         SD1_SB_inst_SD1_SB_bit_inst_58_n111,
         SD1_SB_inst_SD1_SB_bit_inst_58_n110,
         SD1_SB_inst_SD1_SB_bit_inst_58_n109,
         SD1_SB_inst_SD1_SB_bit_inst_58_n108,
         SD1_SB_inst_SD1_SB_bit_inst_58_n107,
         SD1_SB_inst_SD1_SB_bit_inst_58_n106,
         SD1_SB_inst_SD1_SB_bit_inst_58_n105,
         SD1_SB_inst_SD1_SB_bit_inst_58_n104,
         SD1_SB_inst_SD1_SB_bit_inst_58_n103,
         SD1_SB_inst_SD1_SB_bit_inst_58_n102,
         SD1_SB_inst_SD1_SB_bit_inst_58_n101,
         SD1_SB_inst_SD1_SB_bit_inst_58_n100,
         SD1_SB_inst_SD1_SB_bit_inst_58_n99,
         SD1_SB_inst_SD1_SB_bit_inst_58_n98,
         SD1_SB_inst_SD1_SB_bit_inst_58_n97,
         SD1_SB_inst_SD1_SB_bit_inst_59_n141,
         SD1_SB_inst_SD1_SB_bit_inst_59_n140,
         SD1_SB_inst_SD1_SB_bit_inst_59_n139,
         SD1_SB_inst_SD1_SB_bit_inst_59_n138,
         SD1_SB_inst_SD1_SB_bit_inst_59_n137,
         SD1_SB_inst_SD1_SB_bit_inst_59_n136,
         SD1_SB_inst_SD1_SB_bit_inst_59_n135,
         SD1_SB_inst_SD1_SB_bit_inst_59_n134,
         SD1_SB_inst_SD1_SB_bit_inst_59_n133,
         SD1_SB_inst_SD1_SB_bit_inst_59_n132,
         SD1_SB_inst_SD1_SB_bit_inst_59_n131,
         SD1_SB_inst_SD1_SB_bit_inst_59_n130,
         SD1_SB_inst_SD1_SB_bit_inst_59_n129,
         SD1_SB_inst_SD1_SB_bit_inst_59_n128,
         SD1_SB_inst_SD1_SB_bit_inst_59_n127,
         SD1_SB_inst_SD1_SB_bit_inst_59_n126,
         SD1_SB_inst_SD1_SB_bit_inst_59_n125,
         SD1_SB_inst_SD1_SB_bit_inst_59_n124,
         SD1_SB_inst_SD1_SB_bit_inst_59_n123,
         SD1_SB_inst_SD1_SB_bit_inst_59_n122,
         SD1_SB_inst_SD1_SB_bit_inst_59_n121,
         SD1_SB_inst_SD1_SB_bit_inst_59_n120,
         SD1_SB_inst_SD1_SB_bit_inst_59_n119,
         SD1_SB_inst_SD1_SB_bit_inst_59_n118,
         SD1_SB_inst_SD1_SB_bit_inst_59_n117,
         SD1_SB_inst_SD1_SB_bit_inst_59_n116,
         SD1_SB_inst_SD1_SB_bit_inst_59_n115,
         SD1_SB_inst_SD1_SB_bit_inst_59_n114,
         SD1_SB_inst_SD1_SB_bit_inst_59_n113,
         SD1_SB_inst_SD1_SB_bit_inst_59_n112,
         SD1_SB_inst_SD1_SB_bit_inst_59_n111,
         SD1_SB_inst_SD1_SB_bit_inst_59_n110,
         SD1_SB_inst_SD1_SB_bit_inst_59_n109,
         SD1_SB_inst_SD1_SB_bit_inst_59_n108,
         SD1_SB_inst_SD1_SB_bit_inst_59_n107,
         SD1_SB_inst_SD1_SB_bit_inst_59_n106,
         SD1_SB_inst_SD1_SB_bit_inst_59_n105,
         SD1_SB_inst_SD1_SB_bit_inst_59_n104,
         SD1_SB_inst_SD1_SB_bit_inst_59_n103,
         SD1_SB_inst_SD1_SB_bit_inst_59_n102,
         SD1_SB_inst_SD1_SB_bit_inst_59_n101,
         SD1_SB_inst_SD1_SB_bit_inst_59_n100,
         SD1_SB_inst_SD1_SB_bit_inst_60_n131,
         SD1_SB_inst_SD1_SB_bit_inst_60_n130,
         SD1_SB_inst_SD1_SB_bit_inst_60_n129,
         SD1_SB_inst_SD1_SB_bit_inst_60_n128,
         SD1_SB_inst_SD1_SB_bit_inst_60_n127,
         SD1_SB_inst_SD1_SB_bit_inst_60_n126,
         SD1_SB_inst_SD1_SB_bit_inst_60_n125,
         SD1_SB_inst_SD1_SB_bit_inst_60_n124,
         SD1_SB_inst_SD1_SB_bit_inst_60_n123,
         SD1_SB_inst_SD1_SB_bit_inst_60_n122,
         SD1_SB_inst_SD1_SB_bit_inst_60_n121,
         SD1_SB_inst_SD1_SB_bit_inst_60_n120,
         SD1_SB_inst_SD1_SB_bit_inst_60_n119,
         SD1_SB_inst_SD1_SB_bit_inst_60_n118,
         SD1_SB_inst_SD1_SB_bit_inst_60_n117,
         SD1_SB_inst_SD1_SB_bit_inst_60_n116,
         SD1_SB_inst_SD1_SB_bit_inst_60_n115,
         SD1_SB_inst_SD1_SB_bit_inst_60_n114,
         SD1_SB_inst_SD1_SB_bit_inst_60_n113,
         SD1_SB_inst_SD1_SB_bit_inst_60_n112,
         SD1_SB_inst_SD1_SB_bit_inst_60_n111,
         SD1_SB_inst_SD1_SB_bit_inst_60_n110,
         SD1_SB_inst_SD1_SB_bit_inst_60_n109,
         SD1_SB_inst_SD1_SB_bit_inst_60_n108,
         SD1_SB_inst_SD1_SB_bit_inst_60_n107,
         SD1_SB_inst_SD1_SB_bit_inst_60_n106,
         SD1_SB_inst_SD1_SB_bit_inst_60_n105,
         SD1_SB_inst_SD1_SB_bit_inst_60_n104,
         SD1_SB_inst_SD1_SB_bit_inst_60_n103,
         SD1_SB_inst_SD1_SB_bit_inst_60_n102,
         SD1_SB_inst_SD1_SB_bit_inst_60_n101,
         SD1_SB_inst_SD1_SB_bit_inst_60_n100,
         SD1_SB_inst_SD1_SB_bit_inst_60_n99,
         SD1_SB_inst_SD1_SB_bit_inst_60_n98,
         SD1_SB_inst_SD1_SB_bit_inst_60_n97,
         SD1_SB_inst_SD1_SB_bit_inst_60_n96,
         SD1_SB_inst_SD1_SB_bit_inst_60_n95,
         SD1_SB_inst_SD1_SB_bit_inst_60_n94,
         SD1_SB_inst_SD1_SB_bit_inst_60_n93,
         SD1_SB_inst_SD1_SB_bit_inst_60_n92,
         SD1_SB_inst_SD1_SB_bit_inst_61_n110,
         SD1_SB_inst_SD1_SB_bit_inst_61_n109,
         SD1_SB_inst_SD1_SB_bit_inst_61_n108,
         SD1_SB_inst_SD1_SB_bit_inst_61_n107,
         SD1_SB_inst_SD1_SB_bit_inst_61_n106,
         SD1_SB_inst_SD1_SB_bit_inst_61_n105,
         SD1_SB_inst_SD1_SB_bit_inst_61_n104,
         SD1_SB_inst_SD1_SB_bit_inst_61_n103,
         SD1_SB_inst_SD1_SB_bit_inst_61_n102,
         SD1_SB_inst_SD1_SB_bit_inst_61_n101,
         SD1_SB_inst_SD1_SB_bit_inst_61_n100,
         SD1_SB_inst_SD1_SB_bit_inst_61_n99,
         SD1_SB_inst_SD1_SB_bit_inst_61_n98,
         SD1_SB_inst_SD1_SB_bit_inst_61_n97,
         SD1_SB_inst_SD1_SB_bit_inst_61_n96,
         SD1_SB_inst_SD1_SB_bit_inst_61_n95,
         SD1_SB_inst_SD1_SB_bit_inst_61_n94,
         SD1_SB_inst_SD1_SB_bit_inst_61_n93,
         SD1_SB_inst_SD1_SB_bit_inst_61_n92,
         SD1_SB_inst_SD1_SB_bit_inst_61_n91,
         SD1_SB_inst_SD1_SB_bit_inst_61_n90,
         SD1_SB_inst_SD1_SB_bit_inst_61_n89,
         SD1_SB_inst_SD1_SB_bit_inst_61_n88,
         SD1_SB_inst_SD1_SB_bit_inst_61_n87,
         SD1_SB_inst_SD1_SB_bit_inst_61_n86,
         SD1_SB_inst_SD1_SB_bit_inst_61_n85,
         SD1_SB_inst_SD1_SB_bit_inst_61_n84,
         SD1_SB_inst_SD1_SB_bit_inst_61_n83,
         SD1_SB_inst_SD1_SB_bit_inst_61_n82,
         SD1_SB_inst_SD1_SB_bit_inst_61_n81,
         SD1_SB_inst_SD1_SB_bit_inst_61_n80,
         SD1_SB_inst_SD1_SB_bit_inst_61_n79,
         SD1_SB_inst_SD1_SB_bit_inst_61_n78,
         SD1_SB_inst_SD1_SB_bit_inst_61_n77,
         SD1_SB_inst_SD1_SB_bit_inst_62_n138,
         SD1_SB_inst_SD1_SB_bit_inst_62_n137,
         SD1_SB_inst_SD1_SB_bit_inst_62_n136,
         SD1_SB_inst_SD1_SB_bit_inst_62_n135,
         SD1_SB_inst_SD1_SB_bit_inst_62_n134,
         SD1_SB_inst_SD1_SB_bit_inst_62_n133,
         SD1_SB_inst_SD1_SB_bit_inst_62_n132,
         SD1_SB_inst_SD1_SB_bit_inst_62_n131,
         SD1_SB_inst_SD1_SB_bit_inst_62_n130,
         SD1_SB_inst_SD1_SB_bit_inst_62_n129,
         SD1_SB_inst_SD1_SB_bit_inst_62_n128,
         SD1_SB_inst_SD1_SB_bit_inst_62_n127,
         SD1_SB_inst_SD1_SB_bit_inst_62_n126,
         SD1_SB_inst_SD1_SB_bit_inst_62_n125,
         SD1_SB_inst_SD1_SB_bit_inst_62_n124,
         SD1_SB_inst_SD1_SB_bit_inst_62_n123,
         SD1_SB_inst_SD1_SB_bit_inst_62_n122,
         SD1_SB_inst_SD1_SB_bit_inst_62_n121,
         SD1_SB_inst_SD1_SB_bit_inst_62_n120,
         SD1_SB_inst_SD1_SB_bit_inst_62_n119,
         SD1_SB_inst_SD1_SB_bit_inst_62_n118,
         SD1_SB_inst_SD1_SB_bit_inst_62_n117,
         SD1_SB_inst_SD1_SB_bit_inst_62_n116,
         SD1_SB_inst_SD1_SB_bit_inst_62_n115,
         SD1_SB_inst_SD1_SB_bit_inst_62_n114,
         SD1_SB_inst_SD1_SB_bit_inst_62_n113,
         SD1_SB_inst_SD1_SB_bit_inst_62_n112,
         SD1_SB_inst_SD1_SB_bit_inst_62_n111,
         SD1_SB_inst_SD1_SB_bit_inst_62_n110,
         SD1_SB_inst_SD1_SB_bit_inst_62_n109,
         SD1_SB_inst_SD1_SB_bit_inst_62_n108,
         SD1_SB_inst_SD1_SB_bit_inst_62_n107,
         SD1_SB_inst_SD1_SB_bit_inst_62_n106,
         SD1_SB_inst_SD1_SB_bit_inst_62_n105,
         SD1_SB_inst_SD1_SB_bit_inst_62_n104,
         SD1_SB_inst_SD1_SB_bit_inst_62_n103,
         SD1_SB_inst_SD1_SB_bit_inst_62_n102,
         SD1_SB_inst_SD1_SB_bit_inst_62_n101,
         SD1_SB_inst_SD1_SB_bit_inst_62_n100,
         SD1_SB_inst_SD1_SB_bit_inst_62_n99,
         SD1_SB_inst_SD1_SB_bit_inst_62_n98,
         SD1_SB_inst_SD1_SB_bit_inst_62_n97,
         SD1_SB_inst_SD1_SB_bit_inst_63_n141,
         SD1_SB_inst_SD1_SB_bit_inst_63_n140,
         SD1_SB_inst_SD1_SB_bit_inst_63_n139,
         SD1_SB_inst_SD1_SB_bit_inst_63_n138,
         SD1_SB_inst_SD1_SB_bit_inst_63_n137,
         SD1_SB_inst_SD1_SB_bit_inst_63_n136,
         SD1_SB_inst_SD1_SB_bit_inst_63_n135,
         SD1_SB_inst_SD1_SB_bit_inst_63_n134,
         SD1_SB_inst_SD1_SB_bit_inst_63_n133,
         SD1_SB_inst_SD1_SB_bit_inst_63_n132,
         SD1_SB_inst_SD1_SB_bit_inst_63_n131,
         SD1_SB_inst_SD1_SB_bit_inst_63_n130,
         SD1_SB_inst_SD1_SB_bit_inst_63_n129,
         SD1_SB_inst_SD1_SB_bit_inst_63_n128,
         SD1_SB_inst_SD1_SB_bit_inst_63_n127,
         SD1_SB_inst_SD1_SB_bit_inst_63_n126,
         SD1_SB_inst_SD1_SB_bit_inst_63_n125,
         SD1_SB_inst_SD1_SB_bit_inst_63_n124,
         SD1_SB_inst_SD1_SB_bit_inst_63_n123,
         SD1_SB_inst_SD1_SB_bit_inst_63_n122,
         SD1_SB_inst_SD1_SB_bit_inst_63_n121,
         SD1_SB_inst_SD1_SB_bit_inst_63_n120,
         SD1_SB_inst_SD1_SB_bit_inst_63_n119,
         SD1_SB_inst_SD1_SB_bit_inst_63_n118,
         SD1_SB_inst_SD1_SB_bit_inst_63_n117,
         SD1_SB_inst_SD1_SB_bit_inst_63_n116,
         SD1_SB_inst_SD1_SB_bit_inst_63_n115,
         SD1_SB_inst_SD1_SB_bit_inst_63_n114,
         SD1_SB_inst_SD1_SB_bit_inst_63_n113,
         SD1_SB_inst_SD1_SB_bit_inst_63_n112,
         SD1_SB_inst_SD1_SB_bit_inst_63_n111,
         SD1_SB_inst_SD1_SB_bit_inst_63_n110,
         SD1_SB_inst_SD1_SB_bit_inst_63_n109,
         SD1_SB_inst_SD1_SB_bit_inst_63_n108,
         SD1_SB_inst_SD1_SB_bit_inst_63_n107,
         SD1_SB_inst_SD1_SB_bit_inst_63_n106,
         SD1_SB_inst_SD1_SB_bit_inst_63_n105,
         SD1_SB_inst_SD1_SB_bit_inst_63_n104,
         SD1_SB_inst_SD1_SB_bit_inst_63_n103,
         SD1_SB_inst_SD1_SB_bit_inst_63_n102,
         SD1_SB_inst_SD1_SB_bit_inst_63_n101,
         SD1_SB_inst_SD1_SB_bit_inst_63_n100,
         Red_PlaintextInst_LFInst_0_LFInst_0_n3,
         Red_PlaintextInst_LFInst_0_LFInst_1_n3,
         Red_PlaintextInst_LFInst_1_LFInst_0_n3,
         Red_PlaintextInst_LFInst_1_LFInst_1_n3,
         Red_PlaintextInst_LFInst_2_LFInst_0_n3,
         Red_PlaintextInst_LFInst_2_LFInst_1_n3,
         Red_PlaintextInst_LFInst_3_LFInst_0_n3,
         Red_PlaintextInst_LFInst_3_LFInst_1_n3,
         Red_PlaintextInst_LFInst_4_LFInst_0_n3,
         Red_PlaintextInst_LFInst_4_LFInst_1_n3,
         Red_PlaintextInst_LFInst_5_LFInst_0_n3,
         Red_PlaintextInst_LFInst_5_LFInst_1_n3,
         Red_PlaintextInst_LFInst_6_LFInst_0_n3,
         Red_PlaintextInst_LFInst_6_LFInst_1_n3,
         Red_PlaintextInst_LFInst_7_LFInst_0_n3,
         Red_PlaintextInst_LFInst_7_LFInst_1_n3,
         Red_PlaintextInst_LFInst_8_LFInst_0_n3,
         Red_PlaintextInst_LFInst_8_LFInst_1_n3,
         Red_PlaintextInst_LFInst_9_LFInst_0_n3,
         Red_PlaintextInst_LFInst_9_LFInst_1_n3,
         Red_PlaintextInst_LFInst_10_LFInst_0_n3,
         Red_PlaintextInst_LFInst_10_LFInst_1_n3,
         Red_PlaintextInst_LFInst_11_LFInst_0_n3,
         Red_PlaintextInst_LFInst_11_LFInst_1_n3,
         Red_PlaintextInst_LFInst_12_LFInst_0_n3,
         Red_PlaintextInst_LFInst_12_LFInst_1_n3,
         Red_PlaintextInst_LFInst_13_LFInst_0_n3,
         Red_PlaintextInst_LFInst_13_LFInst_1_n3,
         Red_PlaintextInst_LFInst_14_LFInst_0_n3,
         Red_PlaintextInst_LFInst_14_LFInst_1_n3,
         Red_PlaintextInst_LFInst_15_LFInst_0_n3,
         Red_PlaintextInst_LFInst_15_LFInst_1_n3, Red_MCInst_XOR_r0_Inst_0_n5,
         Red_MCInst_XOR_r0_Inst_1_n5, Red_MCInst_XOR_r0_Inst_2_n5,
         Red_MCInst_XOR_r0_Inst_3_n5, Red_MCInst_XOR_r0_Inst_4_n5,
         Red_MCInst_XOR_r0_Inst_5_n5, Red_MCInst_XOR_r0_Inst_6_n5,
         Red_MCInst_XOR_r0_Inst_7_n5, Red_MCInst_XOR_r0_Inst_8_n5,
         Red_MCInst_XOR_r0_Inst_9_n5, Red_MCInst_XOR_r0_Inst_10_n5,
         Red_MCInst_XOR_r0_Inst_11_n5, Red_MCInst_XOR_r0_Inst_12_n5,
         Red_MCInst_XOR_r0_Inst_13_n5, Red_MCInst_XOR_r0_Inst_14_n5,
         Red_MCInst_XOR_r0_Inst_15_n5, Red_MCInst_XOR_r0_Inst_16_n5,
         Red_MCInst_XOR_r0_Inst_17_n5, Red_MCInst_XOR_r0_Inst_18_n5,
         Red_MCInst_XOR_r0_Inst_19_n5, Red_MCInst_XOR_r0_Inst_20_n5,
         Red_MCInst_XOR_r0_Inst_21_n5, Red_MCInst_XOR_r0_Inst_22_n5,
         Red_MCInst_XOR_r0_Inst_23_n5, Red_MCInst_XOR_r0_Inst_24_n5,
         Red_MCInst_XOR_r0_Inst_25_n5, Red_MCInst_XOR_r0_Inst_26_n5,
         Red_MCInst_XOR_r0_Inst_27_n5, Red_AddKeyConstXOR_XORInst_0_0_n5,
         Red_AddKeyConstXOR_XORInst_0_1_n5, Red_AddKeyConstXOR_XORInst_0_2_n5,
         Red_AddKeyConstXOR_XORInst_0_3_n5, Red_AddKeyConstXOR_XORInst_0_4_n5,
         Red_AddKeyConstXOR_XORInst_0_5_n5, Red_AddKeyConstXOR_XORInst_0_6_n5,
         Red_AddKeyConstXOR_XORInst_1_0_n5, Red_AddKeyConstXOR_XORInst_1_1_n5,
         Red_AddKeyConstXOR_XORInst_1_2_n5, Red_AddKeyConstXOR_XORInst_1_3_n5,
         Red_AddKeyConstXOR_XORInst_1_4_n5, Red_AddKeyConstXOR_XORInst_1_5_n5,
         Red_AddKeyConstXOR_XORInst_1_6_n5, F_SD2_RedSB_inst_n80,
         F_SD2_RedSB_inst_n79, F_SD2_RedSB_inst_n78, F_SD2_RedSB_inst_n77,
         F_SD2_RedSB_inst_n76, F_SD2_RedSB_inst_n75, F_SD2_RedSB_inst_n74,
         F_SD2_RedSB_inst_n73, F_SD2_RedSB_inst_n72, F_SD2_RedSB_inst_n71,
         F_SD2_RedSB_inst_n70, F_SD2_RedSB_inst_n69, F_SD2_RedSB_inst_n68,
         F_SD2_RedSB_inst_n67, F_SD2_RedSB_inst_n66, F_SD2_RedSB_inst_n65,
         F_SD2_RedSB_inst_n64, F_SD2_RedSB_inst_n63, F_SD2_RedSB_inst_n62,
         F_SD2_RedSB_inst_n61, F_SD2_RedSB_inst_n60, F_SD2_RedSB_inst_n59,
         F_SD2_RedSB_inst_n58, F_SD2_RedSB_inst_n57, F_SD2_RedSB_inst_n56,
         F_SD2_RedSB_inst_n55, F_SD2_RedSB_inst_n54, F_SD2_RedSB_inst_n53,
         F_SD2_RedSB_inst_n52, F_SD2_RedSB_inst_n51, F_SD2_RedSB_inst_n50,
         F_SD2_RedSB_inst_n49, F_SD2_RedSB_inst_n48, F_SD2_RedSB_inst_n47,
         F_SD2_RedSB_inst_n46, F_SD2_RedSB_inst_n45, F_SD2_RedSB_inst_n44,
         F_SD2_RedSB_inst_n43, F_SD2_RedSB_inst_n42, F_SD2_RedSB_inst_n41,
         F_SD2_RedSB_inst_n40, F_SD2_RedSB_inst_n39, F_SD2_RedSB_inst_n38,
         F_SD2_RedSB_inst_n37, F_SD2_RedSB_inst_n36, F_SD2_RedSB_inst_n35,
         F_SD2_RedSB_inst_n34, F_SD2_RedSB_inst_n33, F_SD2_RedSB_inst_n32,
         F_SD2_RedSB_inst_n31, F_SD2_RedSB_inst_n30, F_SD2_RedSB_inst_n29,
         F_SD2_RedSB_inst_n28, F_SD2_RedSB_inst_n27, F_SD2_RedSB_inst_n26,
         F_SD2_RedSB_inst_n25, F_SD2_RedSB_inst_n24, F_SD2_RedSB_inst_n23,
         F_SD2_RedSB_inst_n22, F_SD2_RedSB_inst_n21, F_SD2_RedSB_inst_n20,
         F_SD2_RedSB_inst_n19, F_SD2_RedSB_inst_n18, F_SD2_RedSB_inst_n17,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n280,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n279,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n278,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n277,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n276,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n275,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n274,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n273,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n272,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n271,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n270,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n269,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n268,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n267,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n266,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n265,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n264,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n263,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n262,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n261,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n260,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n259,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n258,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n257,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n256,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n255,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n254,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n253,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n252,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n251,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n250,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n249,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n248,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n247,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n246,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n245,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n244,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n243,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n242,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n241,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n240,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n239,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n238,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n237,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n236,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n235,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n234,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n233,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n232,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n231,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n230,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n229,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n228,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n227,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n226,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n225,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n224,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n223,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n222,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n221,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n220,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n219,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n218,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n217,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n216,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n215,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n278,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n277,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n276,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n275,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n274,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n273,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n272,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n271,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n270,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n269,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n268,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n267,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n266,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n265,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n264,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n263,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n262,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n261,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n260,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n259,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n258,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n257,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n256,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n255,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n254,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n253,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n252,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n251,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n250,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n249,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n248,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n247,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n246,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n245,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n244,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n243,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n242,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n241,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n240,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n239,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n238,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n237,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n236,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n235,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n234,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n233,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n232,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n231,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n230,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n229,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n228,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n227,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n226,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n225,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n224,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n223,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n222,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n221,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n220,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n219,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n218,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n217,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n216,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n215,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n214,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n240,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n239,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n238,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n237,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n236,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n235,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n234,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n233,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n232,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n231,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n230,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n229,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n228,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n227,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n226,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n225,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n224,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n223,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n222,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n221,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n220,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n219,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n218,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n217,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n216,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n215,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n214,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n213,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n212,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n211,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n210,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n209,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n208,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n207,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n206,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n205,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n204,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n203,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n202,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n201,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n200,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n199,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n198,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n197,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n196,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n195,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n194,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n193,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n192,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n191,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n190,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n290,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n289,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n288,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n287,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n286,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n285,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n284,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n283,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n282,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n281,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n280,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n279,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n278,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n277,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n276,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n275,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n274,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n273,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n272,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n271,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n270,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n269,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n268,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n267,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n266,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n265,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n264,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n263,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n262,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n261,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n260,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n259,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n258,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n257,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n256,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n255,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n254,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n253,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n252,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n251,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n250,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n249,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n248,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n247,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n246,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n245,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n244,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n243,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n242,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n241,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n240,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n239,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n238,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n237,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n236,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n235,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n234,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n233,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n232,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n231,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n230,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n229,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n228,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n227,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n226,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n225,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n224,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n286,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n285,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n284,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n283,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n282,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n281,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n280,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n279,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n278,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n277,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n276,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n275,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n274,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n273,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n272,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n271,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n270,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n269,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n268,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n267,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n266,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n265,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n264,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n263,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n262,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n261,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n260,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n259,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n258,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n257,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n256,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n255,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n254,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n253,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n252,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n251,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n250,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n249,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n248,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n247,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n246,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n245,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n244,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n243,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n242,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n241,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n240,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n239,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n238,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n237,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n236,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n235,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n234,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n233,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n232,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n231,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n230,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n229,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n228,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n227,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n226,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n225,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n224,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n223,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n222,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n221,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n220,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n219,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n218,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n217,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n284,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n283,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n282,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n281,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n280,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n279,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n278,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n277,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n276,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n275,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n274,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n273,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n272,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n271,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n270,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n269,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n268,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n267,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n266,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n265,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n264,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n263,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n262,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n261,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n260,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n259,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n258,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n257,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n256,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n255,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n254,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n253,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n252,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n251,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n250,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n249,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n248,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n247,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n246,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n245,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n244,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n243,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n242,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n241,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n240,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n239,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n238,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n237,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n236,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n235,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n234,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n233,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n232,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n231,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n230,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n229,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n228,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n227,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n226,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n225,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n224,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n223,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n222,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n221,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n220,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n219,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n218,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n217,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n216,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n215,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n176,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n175,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n174,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n173,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n172,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n171,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n170,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n169,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n168,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n167,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n166,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n165,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n164,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n163,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n162,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n161,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n160,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n159,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n158,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n157,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n156,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n155,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n154,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n153,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n152,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n151,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n150,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n149,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n148,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n147,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n146,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n145,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n144,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n143,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n142,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n141,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n140,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n139,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n138,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n137,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n136,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n135,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n134,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n133,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n132,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n131,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n130,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n129,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n128,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n127,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n126,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n125,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n124,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n123,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n122,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n121,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n120,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n119,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n118,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n117,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n116,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n115,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n280,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n279,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n278,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n277,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n276,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n275,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n274,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n273,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n272,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n271,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n270,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n269,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n268,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n267,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n266,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n265,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n264,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n263,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n262,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n261,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n260,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n259,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n258,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n257,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n256,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n255,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n254,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n253,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n252,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n251,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n250,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n249,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n248,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n247,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n246,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n245,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n244,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n243,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n242,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n241,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n240,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n239,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n238,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n237,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n236,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n235,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n234,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n233,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n232,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n231,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n230,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n229,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n228,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n227,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n226,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n225,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n224,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n223,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n222,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n221,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n220,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n219,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n218,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n217,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n216,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n215,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n278,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n277,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n276,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n275,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n274,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n273,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n272,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n271,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n270,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n269,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n268,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n267,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n266,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n265,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n264,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n263,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n262,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n261,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n260,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n259,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n258,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n257,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n256,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n255,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n254,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n253,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n252,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n251,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n250,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n249,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n248,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n247,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n246,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n245,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n244,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n243,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n242,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n241,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n240,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n239,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n238,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n237,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n236,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n235,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n234,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n233,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n232,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n231,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n230,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n229,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n228,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n227,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n226,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n225,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n224,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n223,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n222,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n221,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n220,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n219,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n218,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n217,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n216,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n215,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n214,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n240,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n239,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n238,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n237,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n236,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n235,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n234,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n233,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n232,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n231,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n230,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n229,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n228,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n227,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n226,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n225,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n224,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n223,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n222,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n221,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n220,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n219,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n218,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n217,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n216,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n215,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n214,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n213,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n212,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n211,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n210,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n209,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n208,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n207,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n206,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n205,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n204,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n203,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n202,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n201,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n200,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n199,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n198,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n197,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n196,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n195,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n194,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n193,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n192,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n191,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n190,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n290,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n289,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n288,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n287,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n286,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n285,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n284,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n283,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n282,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n281,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n280,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n279,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n278,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n277,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n276,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n275,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n274,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n273,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n272,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n271,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n270,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n269,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n268,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n267,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n266,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n265,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n264,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n263,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n262,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n261,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n260,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n259,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n258,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n257,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n256,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n255,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n254,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n253,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n252,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n251,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n250,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n249,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n248,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n247,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n246,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n245,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n244,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n243,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n242,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n241,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n240,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n239,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n238,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n237,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n236,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n235,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n234,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n233,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n232,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n231,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n230,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n229,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n228,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n227,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n226,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n225,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n224,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n286,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n285,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n284,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n283,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n282,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n281,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n280,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n279,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n278,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n277,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n276,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n275,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n274,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n273,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n272,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n271,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n270,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n269,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n268,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n267,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n266,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n265,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n264,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n263,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n262,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n261,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n260,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n259,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n258,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n257,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n256,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n255,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n254,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n253,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n252,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n251,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n250,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n249,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n248,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n247,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n246,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n245,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n244,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n243,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n242,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n241,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n240,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n239,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n238,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n237,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n236,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n235,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n234,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n233,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n232,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n231,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n230,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n229,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n228,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n227,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n226,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n225,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n224,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n223,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n222,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n221,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n220,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n219,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n218,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n217,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n284,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n283,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n282,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n281,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n280,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n279,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n278,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n277,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n276,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n275,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n274,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n273,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n272,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n271,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n270,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n269,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n268,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n267,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n266,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n265,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n264,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n263,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n262,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n261,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n260,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n259,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n258,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n257,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n256,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n255,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n254,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n253,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n252,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n251,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n250,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n249,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n248,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n247,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n246,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n245,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n244,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n243,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n242,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n241,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n240,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n239,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n238,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n237,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n236,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n235,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n234,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n233,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n232,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n231,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n230,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n229,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n228,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n227,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n226,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n225,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n224,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n223,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n222,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n221,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n220,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n219,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n218,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n217,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n216,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n215,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n283,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n282,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n281,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n280,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n279,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n278,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n277,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n276,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n275,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n274,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n273,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n272,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n271,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n270,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n269,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n268,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n267,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n266,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n265,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n264,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n263,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n262,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n261,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n260,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n259,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n258,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n257,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n256,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n255,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n254,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n253,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n252,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n251,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n250,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n249,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n248,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n247,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n246,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n245,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n244,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n243,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n242,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n241,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n240,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n239,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n238,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n237,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n236,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n235,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n234,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n233,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n232,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n231,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n230,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n229,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n228,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n227,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n226,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n225,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n224,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n223,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n222,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n280,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n279,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n278,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n277,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n276,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n275,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n274,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n273,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n272,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n271,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n270,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n269,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n268,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n267,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n266,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n265,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n264,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n263,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n262,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n261,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n260,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n259,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n258,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n257,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n256,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n255,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n254,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n253,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n252,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n251,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n250,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n249,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n248,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n247,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n246,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n245,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n244,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n243,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n242,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n241,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n240,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n239,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n238,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n237,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n236,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n235,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n234,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n233,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n232,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n231,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n230,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n229,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n228,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n227,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n226,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n225,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n224,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n223,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n222,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n221,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n220,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n219,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n218,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n217,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n216,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n215,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n278,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n277,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n276,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n275,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n274,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n273,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n272,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n271,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n270,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n269,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n268,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n267,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n266,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n265,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n264,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n263,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n262,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n261,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n260,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n259,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n258,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n257,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n256,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n255,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n254,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n253,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n252,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n251,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n250,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n249,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n248,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n247,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n246,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n245,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n244,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n243,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n242,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n241,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n240,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n239,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n238,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n237,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n236,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n235,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n234,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n233,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n232,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n231,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n230,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n229,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n228,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n227,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n226,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n225,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n224,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n223,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n222,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n221,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n220,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n219,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n218,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n217,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n216,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n215,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n214,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n240,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n239,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n238,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n237,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n236,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n235,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n234,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n233,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n232,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n231,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n230,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n229,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n228,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n227,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n226,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n225,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n224,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n223,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n222,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n221,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n220,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n219,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n218,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n217,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n216,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n215,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n214,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n213,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n212,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n211,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n210,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n209,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n208,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n207,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n206,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n205,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n204,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n203,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n202,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n201,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n200,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n199,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n198,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n197,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n196,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n195,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n194,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n193,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n192,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n191,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n190,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n290,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n289,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n288,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n287,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n286,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n285,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n284,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n283,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n282,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n281,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n280,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n279,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n278,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n277,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n276,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n275,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n274,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n273,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n272,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n271,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n270,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n269,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n268,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n267,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n266,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n265,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n264,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n263,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n262,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n261,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n260,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n259,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n258,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n257,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n256,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n255,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n254,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n253,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n252,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n251,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n250,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n249,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n248,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n247,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n246,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n245,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n244,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n243,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n242,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n241,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n240,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n239,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n238,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n237,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n236,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n235,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n234,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n233,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n232,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n231,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n230,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n229,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n228,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n227,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n226,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n225,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n224,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n286,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n285,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n284,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n283,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n282,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n281,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n280,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n279,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n278,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n277,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n276,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n275,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n274,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n273,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n272,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n271,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n270,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n269,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n268,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n267,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n266,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n265,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n264,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n263,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n262,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n261,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n260,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n259,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n258,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n257,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n256,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n255,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n254,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n253,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n252,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n251,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n250,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n249,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n248,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n247,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n246,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n245,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n244,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n243,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n242,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n241,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n240,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n239,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n238,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n237,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n236,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n235,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n234,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n233,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n232,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n231,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n230,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n229,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n228,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n227,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n226,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n225,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n224,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n223,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n222,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n221,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n220,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n219,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n218,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n217,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n284,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n283,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n282,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n281,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n280,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n279,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n278,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n277,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n276,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n275,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n274,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n273,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n272,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n271,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n270,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n269,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n268,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n267,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n266,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n265,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n264,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n263,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n262,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n261,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n260,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n259,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n258,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n257,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n256,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n255,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n254,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n253,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n252,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n251,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n250,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n249,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n248,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n247,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n246,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n245,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n244,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n243,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n242,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n241,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n240,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n239,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n238,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n237,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n236,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n235,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n234,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n233,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n232,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n231,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n230,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n229,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n228,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n227,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n226,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n225,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n224,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n223,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n222,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n221,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n220,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n219,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n218,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n217,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n216,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n215,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n283,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n282,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n281,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n280,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n279,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n278,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n277,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n276,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n275,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n274,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n273,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n272,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n271,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n270,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n269,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n268,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n267,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n266,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n265,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n264,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n263,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n262,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n261,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n260,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n259,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n258,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n257,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n256,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n255,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n254,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n253,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n252,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n251,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n250,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n249,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n248,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n247,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n246,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n245,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n244,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n243,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n242,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n241,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n240,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n239,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n238,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n237,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n236,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n235,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n234,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n233,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n232,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n231,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n230,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n229,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n228,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n227,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n226,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n225,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n224,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n223,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n222,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n280,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n279,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n278,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n277,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n276,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n275,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n274,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n273,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n272,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n271,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n270,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n269,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n268,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n267,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n266,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n265,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n264,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n263,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n262,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n261,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n260,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n259,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n258,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n257,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n256,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n255,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n254,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n253,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n252,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n251,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n250,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n249,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n248,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n247,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n246,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n245,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n244,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n243,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n242,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n241,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n240,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n239,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n238,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n237,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n236,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n235,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n234,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n233,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n232,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n231,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n230,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n229,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n228,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n227,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n226,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n225,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n224,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n223,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n222,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n221,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n220,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n219,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n218,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n217,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n216,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n215,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n278,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n277,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n276,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n275,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n274,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n273,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n272,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n271,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n270,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n269,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n268,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n267,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n266,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n265,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n264,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n263,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n262,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n261,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n260,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n259,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n258,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n257,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n256,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n255,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n254,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n253,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n252,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n251,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n250,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n249,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n248,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n247,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n246,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n245,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n244,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n243,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n242,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n241,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n240,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n239,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n238,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n237,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n236,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n235,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n234,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n233,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n232,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n231,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n230,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n229,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n228,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n227,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n226,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n225,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n224,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n223,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n222,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n221,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n220,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n219,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n218,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n217,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n216,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n215,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n214,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n240,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n239,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n238,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n237,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n236,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n235,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n234,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n233,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n232,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n231,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n230,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n229,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n228,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n227,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n226,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n225,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n224,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n223,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n222,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n221,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n220,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n219,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n218,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n217,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n216,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n215,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n214,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n213,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n212,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n211,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n210,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n209,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n208,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n207,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n206,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n205,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n204,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n203,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n202,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n201,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n200,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n199,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n198,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n197,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n196,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n195,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n194,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n193,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n192,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n191,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n190,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n290,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n289,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n288,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n287,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n286,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n285,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n284,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n283,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n282,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n281,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n280,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n279,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n278,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n277,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n276,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n275,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n274,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n273,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n272,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n271,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n270,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n269,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n268,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n267,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n266,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n265,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n264,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n263,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n262,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n261,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n260,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n259,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n258,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n257,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n256,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n255,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n254,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n253,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n252,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n251,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n250,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n249,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n248,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n247,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n246,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n245,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n244,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n243,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n242,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n241,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n240,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n239,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n238,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n237,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n236,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n235,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n234,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n233,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n232,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n231,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n230,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n229,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n228,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n227,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n226,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n225,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n224,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n286,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n285,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n284,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n283,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n282,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n281,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n280,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n279,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n278,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n277,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n276,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n275,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n274,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n273,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n272,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n271,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n270,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n269,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n268,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n267,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n266,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n265,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n264,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n263,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n262,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n261,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n260,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n259,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n258,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n257,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n256,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n255,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n254,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n253,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n252,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n251,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n250,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n249,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n248,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n247,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n246,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n245,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n244,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n243,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n242,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n241,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n240,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n239,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n238,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n237,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n236,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n235,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n234,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n233,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n232,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n231,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n230,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n229,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n228,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n227,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n226,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n225,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n224,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n223,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n222,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n221,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n220,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n219,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n218,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n217,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n284,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n283,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n282,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n281,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n280,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n279,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n278,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n277,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n276,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n275,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n274,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n273,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n272,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n271,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n270,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n269,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n268,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n267,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n266,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n265,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n264,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n263,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n262,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n261,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n260,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n259,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n258,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n257,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n256,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n255,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n254,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n253,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n252,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n251,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n250,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n249,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n248,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n247,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n246,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n245,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n244,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n243,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n242,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n241,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n240,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n239,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n238,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n237,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n236,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n235,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n234,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n233,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n232,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n231,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n230,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n229,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n228,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n227,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n226,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n225,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n224,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n223,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n222,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n221,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n220,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n219,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n218,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n217,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n216,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n215,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n283,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n282,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n281,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n280,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n279,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n278,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n277,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n276,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n275,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n274,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n273,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n272,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n271,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n270,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n269,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n268,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n267,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n266,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n265,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n264,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n263,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n262,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n261,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n260,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n259,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n258,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n257,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n256,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n255,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n254,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n253,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n252,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n251,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n250,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n249,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n248,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n247,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n246,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n245,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n244,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n243,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n242,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n241,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n240,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n239,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n238,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n237,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n236,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n235,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n234,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n233,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n232,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n231,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n230,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n229,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n228,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n227,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n226,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n225,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n224,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n223,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n222,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n280,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n279,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n278,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n277,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n276,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n275,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n274,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n273,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n272,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n271,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n270,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n269,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n268,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n267,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n266,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n265,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n264,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n263,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n262,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n261,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n260,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n259,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n258,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n257,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n256,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n255,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n254,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n253,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n252,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n251,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n250,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n249,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n248,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n247,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n246,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n245,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n244,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n243,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n242,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n241,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n240,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n239,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n238,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n237,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n236,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n235,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n234,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n233,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n232,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n231,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n230,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n229,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n228,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n227,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n226,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n225,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n224,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n223,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n222,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n221,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n220,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n219,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n218,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n217,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n216,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n215,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n277,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n276,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n275,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n274,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n273,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n272,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n271,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n270,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n269,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n268,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n267,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n266,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n265,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n264,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n263,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n262,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n261,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n260,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n259,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n258,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n257,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n256,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n255,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n254,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n253,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n252,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n251,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n250,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n249,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n248,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n247,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n246,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n245,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n244,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n243,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n242,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n241,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n240,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n239,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n238,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n237,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n236,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n235,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n234,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n233,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n232,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n231,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n230,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n229,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n228,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n227,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n226,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n225,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n224,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n223,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n222,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n221,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n220,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n219,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n218,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n217,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n216,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n215,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n214,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n240,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n239,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n238,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n237,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n236,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n235,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n234,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n233,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n232,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n231,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n230,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n229,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n228,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n227,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n226,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n225,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n224,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n223,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n222,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n221,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n220,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n219,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n218,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n217,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n216,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n215,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n214,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n213,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n212,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n211,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n210,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n209,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n208,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n207,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n206,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n205,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n204,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n203,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n202,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n201,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n200,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n199,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n198,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n197,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n196,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n195,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n194,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n193,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n192,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n191,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n190,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n291,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n290,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n289,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n288,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n287,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n286,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n285,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n284,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n283,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n282,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n281,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n280,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n279,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n278,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n277,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n276,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n275,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n274,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n273,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n272,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n271,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n270,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n269,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n268,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n267,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n266,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n265,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n264,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n263,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n262,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n261,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n260,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n259,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n258,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n257,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n256,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n255,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n254,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n253,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n252,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n251,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n250,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n249,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n248,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n247,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n246,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n245,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n244,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n243,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n242,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n241,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n240,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n239,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n238,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n237,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n236,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n235,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n234,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n233,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n232,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n231,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n230,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n229,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n228,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n227,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n226,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n225,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n224,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n287,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n286,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n285,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n284,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n283,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n282,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n281,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n280,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n279,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n278,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n277,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n276,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n275,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n274,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n273,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n272,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n271,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n270,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n269,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n268,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n267,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n266,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n265,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n264,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n263,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n262,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n261,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n260,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n259,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n258,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n257,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n256,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n255,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n254,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n253,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n252,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n251,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n250,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n249,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n248,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n247,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n246,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n245,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n244,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n243,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n242,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n241,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n240,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n239,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n238,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n237,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n236,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n235,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n234,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n233,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n232,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n231,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n230,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n229,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n228,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n227,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n226,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n225,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n224,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n223,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n222,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n221,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n220,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n219,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n218,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n217,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n284,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n283,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n282,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n281,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n280,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n279,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n278,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n277,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n276,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n275,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n274,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n273,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n272,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n271,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n270,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n269,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n268,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n267,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n266,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n265,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n264,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n263,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n262,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n261,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n260,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n259,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n258,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n257,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n256,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n255,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n254,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n253,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n252,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n251,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n250,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n249,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n248,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n247,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n246,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n245,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n244,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n243,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n242,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n241,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n240,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n239,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n238,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n237,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n236,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n235,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n234,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n233,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n232,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n231,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n230,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n229,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n228,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n227,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n226,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n225,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n224,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n223,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n222,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n221,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n220,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n219,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n218,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n217,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n216,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n215,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n283,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n282,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n281,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n280,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n279,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n278,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n277,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n276,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n275,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n274,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n273,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n272,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n271,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n270,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n269,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n268,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n267,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n266,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n265,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n264,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n263,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n262,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n261,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n260,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n259,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n258,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n257,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n256,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n255,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n254,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n253,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n252,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n251,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n250,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n249,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n248,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n247,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n246,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n245,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n244,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n243,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n242,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n241,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n240,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n239,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n238,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n237,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n236,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n235,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n234,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n233,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n232,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n231,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n230,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n229,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n228,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n227,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n226,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n225,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n224,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n223,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n222,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n280,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n279,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n278,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n277,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n276,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n275,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n274,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n273,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n272,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n271,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n270,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n269,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n268,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n267,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n266,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n265,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n264,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n263,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n262,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n261,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n260,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n259,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n258,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n257,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n256,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n255,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n254,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n253,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n252,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n251,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n250,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n249,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n248,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n247,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n246,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n245,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n244,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n243,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n242,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n241,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n240,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n239,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n238,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n237,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n236,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n235,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n234,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n233,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n232,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n231,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n230,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n229,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n228,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n227,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n226,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n225,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n224,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n223,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n222,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n221,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n220,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n219,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n218,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n217,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n216,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n215,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n278,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n277,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n276,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n275,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n274,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n273,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n272,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n271,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n270,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n269,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n268,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n267,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n266,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n265,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n264,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n263,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n262,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n261,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n260,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n259,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n258,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n257,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n256,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n255,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n254,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n253,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n252,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n251,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n250,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n249,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n248,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n247,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n246,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n245,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n244,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n243,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n242,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n241,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n240,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n239,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n238,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n237,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n236,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n235,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n234,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n233,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n232,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n231,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n230,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n229,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n228,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n227,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n226,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n225,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n224,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n223,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n222,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n221,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n220,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n219,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n218,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n217,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n216,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n215,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n214,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n240,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n239,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n238,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n237,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n236,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n235,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n234,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n233,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n232,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n231,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n230,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n229,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n228,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n227,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n226,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n225,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n224,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n223,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n222,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n221,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n220,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n219,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n218,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n217,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n216,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n215,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n214,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n213,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n212,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n211,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n210,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n209,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n208,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n207,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n206,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n205,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n204,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n203,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n202,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n201,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n200,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n199,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n198,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n197,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n196,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n195,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n194,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n193,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n192,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n191,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n190,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n289,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n288,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n287,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n286,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n285,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n284,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n283,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n282,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n281,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n280,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n279,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n278,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n277,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n276,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n275,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n274,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n273,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n272,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n271,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n270,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n269,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n268,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n267,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n266,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n265,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n264,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n263,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n262,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n261,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n260,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n259,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n258,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n257,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n256,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n255,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n254,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n253,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n252,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n251,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n250,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n249,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n248,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n247,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n246,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n245,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n244,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n243,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n242,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n241,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n240,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n239,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n238,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n237,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n236,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n235,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n234,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n233,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n232,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n231,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n230,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n229,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n228,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n227,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n226,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n225,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n224,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n286,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n285,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n284,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n283,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n282,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n281,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n280,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n279,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n278,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n277,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n276,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n275,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n274,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n273,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n272,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n271,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n270,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n269,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n268,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n267,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n266,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n265,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n264,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n263,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n262,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n261,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n260,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n259,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n258,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n257,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n256,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n255,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n254,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n253,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n252,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n251,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n250,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n249,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n248,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n247,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n246,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n245,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n244,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n243,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n242,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n241,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n240,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n239,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n238,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n237,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n236,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n235,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n234,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n233,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n232,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n231,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n230,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n229,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n228,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n227,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n226,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n225,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n224,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n223,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n222,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n221,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n220,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n219,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n218,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n217,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n284,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n283,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n282,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n281,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n280,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n279,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n278,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n277,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n276,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n275,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n274,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n273,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n272,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n271,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n270,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n269,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n268,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n267,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n266,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n265,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n264,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n263,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n262,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n261,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n260,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n259,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n258,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n257,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n256,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n255,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n254,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n253,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n252,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n251,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n250,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n249,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n248,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n247,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n246,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n245,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n244,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n243,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n242,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n241,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n240,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n239,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n238,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n237,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n236,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n235,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n234,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n233,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n232,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n231,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n230,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n229,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n228,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n227,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n226,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n225,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n224,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n223,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n222,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n221,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n220,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n219,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n218,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n217,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n216,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n215,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n283,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n282,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n281,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n280,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n279,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n278,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n277,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n276,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n275,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n274,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n273,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n272,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n271,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n270,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n269,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n268,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n267,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n266,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n265,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n264,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n263,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n262,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n261,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n260,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n259,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n258,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n257,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n256,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n255,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n254,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n253,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n252,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n251,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n250,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n249,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n248,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n247,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n246,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n245,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n244,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n243,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n242,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n241,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n240,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n239,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n238,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n237,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n236,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n235,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n234,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n233,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n232,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n231,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n230,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n229,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n228,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n227,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n226,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n225,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n224,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n223,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n222,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n280,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n279,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n278,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n277,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n276,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n275,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n274,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n273,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n272,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n271,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n270,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n269,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n268,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n267,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n266,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n265,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n264,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n263,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n262,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n261,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n260,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n259,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n258,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n257,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n256,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n255,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n254,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n253,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n252,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n251,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n250,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n249,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n248,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n247,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n246,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n245,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n244,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n243,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n242,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n241,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n240,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n239,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n238,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n237,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n236,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n235,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n234,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n233,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n232,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n231,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n230,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n229,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n228,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n227,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n226,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n225,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n224,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n223,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n222,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n221,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n220,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n219,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n218,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n217,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n216,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n215,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n278,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n277,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n276,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n275,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n274,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n273,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n272,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n271,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n270,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n269,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n268,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n267,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n266,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n265,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n264,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n263,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n262,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n261,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n260,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n259,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n258,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n257,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n256,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n255,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n254,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n253,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n252,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n251,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n250,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n249,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n248,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n247,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n246,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n245,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n244,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n243,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n242,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n241,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n240,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n239,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n238,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n237,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n236,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n235,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n234,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n233,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n232,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n231,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n230,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n229,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n228,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n227,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n226,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n225,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n224,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n223,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n222,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n221,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n220,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n219,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n218,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n217,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n216,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n215,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n214,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n240,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n239,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n238,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n237,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n236,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n235,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n234,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n233,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n232,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n231,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n230,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n229,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n228,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n227,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n226,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n225,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n224,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n223,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n222,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n221,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n220,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n219,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n218,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n217,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n216,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n215,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n214,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n213,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n212,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n211,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n210,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n209,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n208,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n207,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n206,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n205,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n204,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n203,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n202,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n201,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n200,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n199,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n198,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n197,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n196,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n195,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n194,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n193,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n192,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n191,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n190,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n289,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n288,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n287,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n286,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n285,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n284,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n283,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n282,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n281,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n280,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n279,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n278,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n277,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n276,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n275,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n274,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n273,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n272,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n271,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n270,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n269,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n268,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n267,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n266,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n265,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n264,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n263,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n262,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n261,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n260,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n259,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n258,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n257,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n256,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n255,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n254,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n253,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n252,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n251,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n250,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n249,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n248,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n247,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n246,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n245,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n244,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n243,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n242,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n241,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n240,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n239,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n238,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n237,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n236,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n235,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n234,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n233,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n232,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n231,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n230,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n229,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n228,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n227,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n226,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n225,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n224,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n286,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n285,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n284,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n283,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n282,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n281,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n280,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n279,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n278,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n277,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n276,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n275,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n274,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n273,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n272,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n271,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n270,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n269,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n268,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n267,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n266,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n265,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n264,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n263,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n262,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n261,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n260,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n259,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n258,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n257,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n256,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n255,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n254,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n253,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n252,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n251,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n250,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n249,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n248,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n247,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n246,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n245,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n244,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n243,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n242,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n241,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n240,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n239,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n238,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n237,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n236,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n235,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n234,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n233,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n232,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n231,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n230,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n229,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n228,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n227,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n226,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n225,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n224,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n223,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n222,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n221,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n220,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n219,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n218,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n217,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n284,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n283,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n282,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n281,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n280,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n279,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n278,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n277,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n276,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n275,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n274,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n273,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n272,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n271,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n270,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n269,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n268,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n267,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n266,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n265,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n264,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n263,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n262,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n261,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n260,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n259,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n258,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n257,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n256,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n255,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n254,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n253,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n252,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n251,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n250,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n249,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n248,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n247,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n246,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n245,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n244,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n243,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n242,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n241,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n240,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n239,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n238,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n237,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n236,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n235,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n234,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n233,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n232,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n231,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n230,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n229,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n228,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n227,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n226,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n225,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n224,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n223,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n222,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n221,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n220,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n219,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n218,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n217,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n216,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n215,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n283,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n282,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n281,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n280,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n279,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n278,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n277,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n276,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n275,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n274,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n273,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n272,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n271,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n270,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n269,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n268,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n267,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n266,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n265,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n264,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n263,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n262,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n261,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n260,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n259,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n258,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n257,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n256,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n255,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n254,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n253,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n252,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n251,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n250,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n249,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n248,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n247,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n246,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n245,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n244,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n243,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n242,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n241,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n240,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n239,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n238,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n237,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n236,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n235,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n234,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n233,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n232,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n231,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n230,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n229,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n228,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n227,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n226,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n225,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n224,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n223,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n222,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n280,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n279,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n278,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n277,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n276,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n275,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n274,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n273,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n272,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n271,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n270,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n269,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n268,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n267,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n266,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n265,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n264,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n263,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n262,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n261,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n260,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n259,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n258,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n257,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n256,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n255,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n254,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n253,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n252,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n251,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n250,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n249,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n248,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n247,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n246,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n245,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n244,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n243,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n242,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n241,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n240,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n239,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n238,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n237,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n236,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n235,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n234,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n233,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n232,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n231,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n230,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n229,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n228,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n227,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n226,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n225,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n224,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n223,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n222,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n221,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n220,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n219,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n218,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n217,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n216,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n215,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n277,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n276,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n275,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n274,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n273,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n272,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n271,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n270,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n269,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n268,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n267,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n266,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n265,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n264,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n263,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n262,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n261,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n260,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n259,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n258,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n257,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n256,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n255,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n254,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n253,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n252,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n251,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n250,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n249,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n248,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n247,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n246,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n245,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n244,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n243,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n242,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n241,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n240,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n239,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n238,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n237,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n236,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n235,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n234,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n233,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n232,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n231,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n230,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n229,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n228,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n227,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n226,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n225,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n224,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n223,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n222,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n221,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n220,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n219,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n218,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n217,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n216,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n215,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n214,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n240,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n239,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n238,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n237,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n236,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n235,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n234,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n233,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n232,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n231,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n230,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n229,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n228,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n227,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n226,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n225,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n224,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n223,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n222,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n221,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n220,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n219,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n218,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n217,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n216,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n215,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n214,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n213,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n212,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n211,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n210,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n209,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n208,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n207,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n206,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n205,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n204,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n203,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n202,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n201,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n200,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n199,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n198,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n197,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n196,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n195,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n194,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n193,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n192,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n191,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n190,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n291,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n290,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n289,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n288,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n287,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n286,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n285,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n284,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n283,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n282,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n281,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n280,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n279,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n278,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n277,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n276,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n275,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n274,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n273,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n272,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n271,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n270,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n269,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n268,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n267,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n266,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n265,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n264,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n263,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n262,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n261,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n260,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n259,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n258,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n257,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n256,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n255,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n254,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n253,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n252,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n251,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n250,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n249,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n248,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n247,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n246,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n245,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n244,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n243,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n242,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n241,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n240,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n239,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n238,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n237,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n236,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n235,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n234,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n233,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n232,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n231,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n230,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n229,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n228,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n227,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n226,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n225,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n224,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n287,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n286,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n285,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n284,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n283,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n282,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n281,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n280,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n279,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n278,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n277,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n276,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n275,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n274,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n273,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n272,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n271,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n270,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n269,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n268,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n267,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n266,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n265,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n264,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n263,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n262,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n261,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n260,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n259,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n258,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n257,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n256,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n255,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n254,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n253,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n252,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n251,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n250,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n249,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n248,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n247,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n246,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n245,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n244,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n243,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n242,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n241,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n240,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n239,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n238,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n237,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n236,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n235,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n234,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n233,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n232,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n231,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n230,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n229,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n228,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n227,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n226,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n225,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n224,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n223,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n222,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n221,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n220,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n219,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n218,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n217,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n284,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n283,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n282,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n281,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n280,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n279,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n278,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n277,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n276,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n275,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n274,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n273,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n272,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n271,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n270,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n269,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n268,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n267,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n266,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n265,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n264,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n263,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n262,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n261,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n260,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n259,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n258,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n257,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n256,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n255,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n254,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n253,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n252,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n251,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n250,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n249,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n248,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n247,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n246,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n245,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n244,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n243,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n242,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n241,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n240,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n239,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n238,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n237,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n236,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n235,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n234,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n233,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n232,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n231,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n230,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n229,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n228,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n227,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n226,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n225,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n224,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n223,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n222,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n221,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n220,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n219,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n218,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n217,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n216,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n215,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n283,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n282,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n281,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n280,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n279,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n278,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n277,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n276,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n275,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n274,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n273,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n272,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n271,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n270,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n269,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n268,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n267,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n266,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n265,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n264,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n263,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n262,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n261,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n260,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n259,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n258,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n257,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n256,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n255,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n254,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n253,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n252,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n251,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n250,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n249,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n248,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n247,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n246,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n245,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n244,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n243,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n242,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n241,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n240,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n239,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n238,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n237,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n236,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n235,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n234,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n233,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n232,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n231,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n230,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n229,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n228,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n227,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n226,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n225,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n224,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n223,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n222,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n280,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n279,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n278,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n277,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n276,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n275,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n274,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n273,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n272,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n271,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n270,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n269,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n268,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n267,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n266,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n265,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n264,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n263,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n262,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n261,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n260,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n259,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n258,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n257,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n256,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n255,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n254,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n253,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n252,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n251,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n250,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n249,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n248,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n247,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n246,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n245,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n244,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n243,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n242,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n241,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n240,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n239,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n238,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n237,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n236,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n235,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n234,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n233,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n232,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n231,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n230,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n229,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n228,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n227,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n226,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n225,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n224,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n223,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n222,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n221,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n220,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n219,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n218,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n217,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n216,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n215,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n279,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n278,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n277,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n276,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n275,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n274,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n273,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n272,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n271,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n270,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n269,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n268,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n267,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n266,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n265,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n264,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n263,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n262,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n261,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n260,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n259,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n258,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n257,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n256,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n255,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n254,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n253,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n252,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n251,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n250,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n249,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n248,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n247,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n246,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n245,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n244,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n243,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n242,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n241,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n240,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n239,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n238,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n237,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n236,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n235,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n234,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n233,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n232,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n231,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n230,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n229,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n228,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n227,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n226,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n225,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n224,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n223,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n222,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n221,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n220,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n219,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n218,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n217,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n216,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n215,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n214,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n240,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n239,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n238,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n237,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n236,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n235,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n234,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n233,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n232,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n231,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n230,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n229,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n228,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n227,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n226,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n225,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n224,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n223,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n222,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n221,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n220,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n219,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n218,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n217,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n216,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n215,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n214,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n213,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n212,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n211,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n210,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n209,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n208,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n207,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n206,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n205,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n204,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n203,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n202,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n201,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n200,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n199,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n198,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n197,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n196,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n195,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n194,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n193,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n192,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n191,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n190,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n291,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n290,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n289,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n288,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n287,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n286,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n285,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n284,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n283,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n282,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n281,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n280,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n279,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n278,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n277,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n276,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n275,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n274,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n273,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n272,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n271,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n270,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n269,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n268,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n267,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n266,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n265,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n264,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n263,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n262,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n261,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n260,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n259,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n258,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n257,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n256,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n255,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n254,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n253,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n252,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n251,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n250,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n249,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n248,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n247,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n246,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n245,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n244,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n243,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n242,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n241,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n240,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n239,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n238,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n237,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n236,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n235,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n234,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n233,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n232,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n231,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n230,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n229,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n228,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n227,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n226,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n225,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n224,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n286,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n285,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n284,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n283,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n282,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n281,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n280,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n279,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n278,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n277,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n276,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n275,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n274,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n273,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n272,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n271,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n270,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n269,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n268,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n267,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n266,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n265,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n264,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n263,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n262,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n261,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n260,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n259,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n258,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n257,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n256,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n255,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n254,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n253,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n252,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n251,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n250,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n249,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n248,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n247,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n246,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n245,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n244,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n243,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n242,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n241,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n240,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n239,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n238,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n237,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n236,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n235,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n234,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n233,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n232,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n231,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n230,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n229,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n228,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n227,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n226,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n225,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n224,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n223,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n222,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n221,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n220,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n219,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n218,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n217,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n284,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n283,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n282,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n281,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n280,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n279,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n278,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n277,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n276,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n275,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n274,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n273,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n272,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n271,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n270,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n269,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n268,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n267,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n266,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n265,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n264,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n263,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n262,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n261,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n260,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n259,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n258,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n257,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n256,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n255,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n254,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n253,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n252,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n251,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n250,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n249,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n248,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n247,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n246,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n245,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n244,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n243,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n242,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n241,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n240,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n239,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n238,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n237,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n236,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n235,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n234,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n233,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n232,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n231,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n230,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n229,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n228,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n227,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n226,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n225,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n224,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n223,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n222,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n221,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n220,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n219,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n218,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n217,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n216,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n215,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n283,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n282,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n281,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n280,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n279,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n278,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n277,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n276,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n275,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n274,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n273,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n272,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n271,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n270,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n269,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n268,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n267,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n266,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n265,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n264,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n263,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n262,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n261,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n260,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n259,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n258,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n257,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n256,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n255,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n254,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n253,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n252,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n251,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n250,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n249,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n248,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n247,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n246,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n245,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n244,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n243,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n242,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n241,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n240,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n239,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n238,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n237,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n236,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n235,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n234,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n233,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n232,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n231,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n230,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n229,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n228,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n227,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n226,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n225,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n224,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n223,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n222,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n280,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n279,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n278,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n277,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n276,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n275,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n274,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n273,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n272,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n271,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n270,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n269,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n268,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n267,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n266,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n265,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n264,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n263,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n262,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n261,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n260,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n259,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n258,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n257,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n256,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n255,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n254,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n253,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n252,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n251,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n250,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n249,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n248,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n247,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n246,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n245,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n244,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n243,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n242,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n241,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n240,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n239,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n238,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n237,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n236,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n235,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n234,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n233,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n232,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n231,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n230,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n229,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n228,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n227,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n226,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n225,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n224,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n223,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n222,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n221,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n220,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n219,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n218,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n217,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n216,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n215,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n279,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n278,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n277,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n276,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n275,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n274,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n273,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n272,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n271,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n270,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n269,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n268,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n267,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n266,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n265,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n264,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n263,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n262,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n261,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n260,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n259,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n258,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n257,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n256,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n255,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n254,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n253,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n252,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n251,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n250,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n249,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n248,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n247,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n246,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n245,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n244,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n243,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n242,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n241,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n240,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n239,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n238,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n237,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n236,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n235,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n234,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n233,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n232,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n231,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n230,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n229,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n228,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n227,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n226,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n225,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n224,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n223,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n222,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n221,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n220,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n219,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n218,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n217,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n216,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n215,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n214,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n240,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n239,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n238,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n237,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n236,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n235,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n234,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n233,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n232,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n231,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n230,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n229,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n228,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n227,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n226,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n225,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n224,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n223,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n222,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n221,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n220,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n219,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n218,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n217,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n216,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n215,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n214,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n213,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n212,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n211,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n210,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n209,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n208,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n207,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n206,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n205,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n204,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n203,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n202,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n201,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n200,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n199,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n198,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n197,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n196,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n195,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n194,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n193,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n192,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n191,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n190,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n291,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n290,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n289,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n288,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n287,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n286,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n285,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n284,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n283,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n282,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n281,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n280,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n279,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n278,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n277,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n276,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n275,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n274,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n273,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n272,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n271,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n270,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n269,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n268,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n267,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n266,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n265,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n264,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n263,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n262,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n261,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n260,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n259,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n258,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n257,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n256,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n255,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n254,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n253,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n252,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n251,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n250,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n249,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n248,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n247,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n246,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n245,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n244,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n243,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n242,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n241,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n240,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n239,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n238,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n237,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n236,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n235,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n234,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n233,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n232,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n231,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n230,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n229,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n228,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n227,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n226,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n225,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n224,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n286,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n285,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n284,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n283,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n282,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n281,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n280,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n279,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n278,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n277,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n276,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n275,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n274,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n273,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n272,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n271,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n270,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n269,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n268,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n267,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n266,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n265,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n264,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n263,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n262,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n261,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n260,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n259,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n258,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n257,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n256,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n255,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n254,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n253,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n252,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n251,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n250,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n249,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n248,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n247,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n246,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n245,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n244,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n243,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n242,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n241,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n240,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n239,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n238,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n237,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n236,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n235,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n234,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n233,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n232,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n231,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n230,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n229,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n228,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n227,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n226,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n225,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n224,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n223,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n222,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n221,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n220,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n219,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n218,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n217,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n284,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n283,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n282,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n281,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n280,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n279,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n278,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n277,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n276,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n275,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n274,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n273,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n272,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n271,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n270,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n269,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n268,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n267,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n266,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n265,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n264,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n263,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n262,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n261,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n260,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n259,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n258,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n257,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n256,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n255,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n254,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n253,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n252,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n251,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n250,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n249,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n248,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n247,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n246,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n245,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n244,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n243,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n242,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n241,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n240,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n239,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n238,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n237,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n236,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n235,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n234,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n233,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n232,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n231,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n230,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n229,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n228,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n227,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n226,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n225,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n224,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n223,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n222,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n221,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n220,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n219,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n218,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n217,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n216,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n215,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n283,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n282,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n281,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n280,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n279,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n278,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n277,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n276,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n275,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n274,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n273,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n272,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n271,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n270,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n269,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n268,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n267,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n266,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n265,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n264,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n263,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n262,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n261,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n260,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n259,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n258,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n257,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n256,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n255,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n254,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n253,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n252,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n251,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n250,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n249,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n248,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n247,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n246,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n245,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n244,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n243,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n242,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n241,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n240,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n239,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n238,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n237,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n236,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n235,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n234,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n233,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n232,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n231,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n230,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n229,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n228,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n227,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n226,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n225,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n224,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n223,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n222,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n280,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n279,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n278,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n277,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n276,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n275,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n274,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n273,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n272,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n271,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n270,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n269,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n268,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n267,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n266,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n265,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n264,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n263,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n262,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n261,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n260,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n259,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n258,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n257,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n256,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n255,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n254,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n253,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n252,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n251,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n250,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n249,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n248,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n247,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n246,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n245,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n244,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n243,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n242,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n241,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n240,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n239,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n238,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n237,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n236,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n235,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n234,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n233,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n232,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n231,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n230,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n229,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n228,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n227,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n226,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n225,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n224,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n223,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n222,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n221,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n220,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n219,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n218,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n217,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n216,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n215,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n279,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n278,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n277,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n276,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n275,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n274,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n273,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n272,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n271,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n270,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n269,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n268,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n267,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n266,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n265,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n264,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n263,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n262,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n261,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n260,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n259,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n258,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n257,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n256,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n255,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n254,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n253,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n252,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n251,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n250,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n249,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n248,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n247,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n246,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n245,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n244,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n243,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n242,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n241,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n240,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n239,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n238,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n237,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n236,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n235,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n234,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n233,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n232,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n231,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n230,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n229,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n228,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n227,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n226,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n225,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n224,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n223,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n222,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n221,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n220,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n219,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n218,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n217,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n216,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n215,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n214,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n240,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n239,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n238,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n237,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n236,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n235,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n234,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n233,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n232,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n231,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n230,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n229,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n228,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n227,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n226,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n225,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n224,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n223,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n222,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n221,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n220,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n219,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n218,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n217,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n216,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n215,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n214,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n213,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n212,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n211,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n210,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n209,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n208,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n207,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n206,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n205,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n204,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n203,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n202,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n201,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n200,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n199,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n198,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n197,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n196,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n195,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n194,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n193,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n192,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n191,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n190,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n291,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n290,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n289,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n288,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n287,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n286,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n285,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n284,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n283,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n282,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n281,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n280,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n279,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n278,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n277,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n276,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n275,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n274,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n273,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n272,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n271,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n270,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n269,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n268,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n267,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n266,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n265,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n264,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n263,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n262,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n261,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n260,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n259,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n258,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n257,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n256,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n255,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n254,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n253,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n252,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n251,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n250,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n249,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n248,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n247,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n246,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n245,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n244,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n243,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n242,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n241,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n240,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n239,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n238,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n237,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n236,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n235,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n234,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n233,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n232,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n231,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n230,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n229,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n228,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n227,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n226,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n225,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n224,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n286,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n285,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n284,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n283,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n282,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n281,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n280,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n279,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n278,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n277,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n276,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n275,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n274,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n273,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n272,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n271,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n270,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n269,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n268,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n267,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n266,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n265,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n264,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n263,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n262,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n261,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n260,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n259,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n258,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n257,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n256,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n255,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n254,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n253,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n252,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n251,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n250,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n249,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n248,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n247,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n246,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n245,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n244,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n243,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n242,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n241,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n240,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n239,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n238,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n237,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n236,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n235,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n234,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n233,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n232,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n231,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n230,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n229,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n228,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n227,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n226,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n225,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n224,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n223,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n222,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n221,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n220,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n219,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n218,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n217,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n284,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n283,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n282,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n281,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n280,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n279,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n278,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n277,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n276,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n275,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n274,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n273,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n272,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n271,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n270,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n269,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n268,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n267,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n266,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n265,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n264,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n263,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n262,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n261,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n260,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n259,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n258,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n257,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n256,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n255,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n254,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n253,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n252,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n251,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n250,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n249,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n248,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n247,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n246,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n245,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n244,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n243,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n242,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n241,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n240,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n239,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n238,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n237,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n236,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n235,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n234,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n233,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n232,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n231,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n230,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n229,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n228,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n227,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n226,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n225,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n224,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n223,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n222,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n221,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n220,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n219,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n218,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n217,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n216,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n215,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n283,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n282,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n281,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n280,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n279,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n278,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n277,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n276,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n275,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n274,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n273,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n272,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n271,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n270,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n269,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n268,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n267,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n266,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n265,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n264,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n263,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n262,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n261,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n260,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n259,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n258,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n257,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n256,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n255,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n254,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n253,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n252,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n251,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n250,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n249,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n248,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n247,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n246,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n245,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n244,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n243,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n242,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n241,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n240,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n239,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n238,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n237,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n236,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n235,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n234,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n233,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n232,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n231,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n230,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n229,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n228,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n227,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n226,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n225,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n224,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n223,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n222,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n280,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n279,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n278,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n277,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n276,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n275,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n274,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n273,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n272,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n271,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n270,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n269,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n268,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n267,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n266,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n265,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n264,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n263,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n262,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n261,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n260,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n259,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n258,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n257,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n256,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n255,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n254,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n253,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n252,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n251,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n250,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n249,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n248,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n247,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n246,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n245,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n244,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n243,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n242,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n241,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n240,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n239,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n238,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n237,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n236,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n235,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n234,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n233,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n232,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n231,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n230,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n229,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n228,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n227,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n226,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n225,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n224,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n223,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n222,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n221,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n220,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n219,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n218,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n217,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n216,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n215,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n279,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n278,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n277,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n276,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n275,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n274,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n273,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n272,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n271,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n270,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n269,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n268,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n267,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n266,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n265,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n264,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n263,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n262,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n261,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n260,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n259,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n258,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n257,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n256,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n255,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n254,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n253,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n252,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n251,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n250,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n249,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n248,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n247,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n246,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n245,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n244,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n243,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n242,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n241,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n240,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n239,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n238,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n237,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n236,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n235,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n234,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n233,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n232,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n231,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n230,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n229,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n228,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n227,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n226,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n225,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n224,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n223,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n222,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n221,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n220,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n219,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n218,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n217,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n216,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n215,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n214,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n240,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n239,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n238,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n237,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n236,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n235,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n234,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n233,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n232,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n231,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n230,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n229,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n228,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n227,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n226,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n225,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n224,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n223,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n222,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n221,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n220,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n219,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n218,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n217,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n216,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n215,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n214,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n213,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n212,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n211,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n210,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n209,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n208,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n207,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n206,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n205,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n204,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n203,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n202,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n201,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n200,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n199,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n198,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n197,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n196,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n195,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n194,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n193,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n192,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n191,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n190,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n291,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n290,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n289,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n288,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n287,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n286,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n285,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n284,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n283,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n282,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n281,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n280,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n279,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n278,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n277,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n276,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n275,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n274,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n273,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n272,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n271,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n270,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n269,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n268,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n267,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n266,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n265,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n264,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n263,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n262,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n261,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n260,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n259,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n258,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n257,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n256,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n255,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n254,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n253,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n252,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n251,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n250,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n249,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n248,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n247,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n246,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n245,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n244,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n243,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n242,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n241,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n240,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n239,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n238,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n237,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n236,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n235,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n234,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n233,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n232,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n231,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n230,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n229,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n228,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n227,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n226,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n225,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n224,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n286,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n285,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n284,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n283,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n282,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n281,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n280,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n279,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n278,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n277,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n276,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n275,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n274,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n273,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n272,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n271,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n270,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n269,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n268,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n267,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n266,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n265,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n264,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n263,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n262,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n261,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n260,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n259,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n258,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n257,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n256,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n255,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n254,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n253,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n252,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n251,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n250,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n249,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n248,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n247,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n246,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n245,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n244,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n243,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n242,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n241,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n240,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n239,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n238,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n237,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n236,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n235,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n234,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n233,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n232,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n231,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n230,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n229,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n228,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n227,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n226,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n225,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n224,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n223,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n222,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n221,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n220,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n219,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n218,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n217,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n284,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n283,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n282,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n281,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n280,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n279,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n278,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n277,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n276,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n275,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n274,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n273,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n272,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n271,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n270,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n269,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n268,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n267,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n266,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n265,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n264,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n263,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n262,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n261,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n260,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n259,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n258,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n257,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n256,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n255,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n254,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n253,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n252,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n251,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n250,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n249,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n248,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n247,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n246,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n245,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n244,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n243,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n242,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n241,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n240,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n239,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n238,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n237,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n236,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n235,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n234,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n233,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n232,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n231,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n230,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n229,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n228,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n227,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n226,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n225,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n224,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n223,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n222,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n221,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n220,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n219,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n218,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n217,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n216,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n215,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n283,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n282,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n281,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n280,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n279,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n278,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n277,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n276,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n275,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n274,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n273,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n272,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n271,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n270,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n269,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n268,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n267,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n266,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n265,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n264,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n263,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n262,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n261,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n260,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n259,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n258,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n257,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n256,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n255,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n254,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n253,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n252,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n251,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n250,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n249,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n248,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n247,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n246,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n245,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n244,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n243,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n242,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n241,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n240,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n239,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n238,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n237,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n236,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n235,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n234,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n233,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n232,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n231,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n230,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n229,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n228,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n227,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n226,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n225,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n224,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n223,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n222,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n280,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n279,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n278,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n277,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n276,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n275,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n274,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n273,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n272,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n271,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n270,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n269,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n268,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n267,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n266,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n265,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n264,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n263,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n262,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n261,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n260,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n259,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n258,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n257,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n256,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n255,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n254,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n253,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n252,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n251,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n250,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n249,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n248,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n247,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n246,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n245,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n244,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n243,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n242,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n241,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n240,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n239,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n238,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n237,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n236,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n235,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n234,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n233,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n232,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n231,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n230,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n229,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n228,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n227,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n226,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n225,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n224,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n223,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n222,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n221,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n220,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n219,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n218,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n217,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n216,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n215,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n279,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n278,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n277,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n276,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n275,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n274,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n273,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n272,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n271,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n270,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n269,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n268,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n267,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n266,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n265,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n264,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n263,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n262,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n261,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n260,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n259,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n258,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n257,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n256,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n255,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n254,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n253,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n252,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n251,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n250,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n249,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n248,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n247,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n246,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n245,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n244,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n243,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n242,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n241,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n240,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n239,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n238,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n237,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n236,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n235,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n234,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n233,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n232,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n231,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n230,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n229,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n228,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n227,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n226,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n225,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n224,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n223,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n222,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n221,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n220,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n219,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n218,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n217,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n216,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n215,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n214,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n240,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n239,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n238,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n237,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n236,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n235,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n234,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n233,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n232,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n231,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n230,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n229,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n228,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n227,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n226,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n225,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n224,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n223,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n222,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n221,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n220,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n219,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n218,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n217,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n216,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n215,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n214,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n213,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n212,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n211,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n210,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n209,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n208,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n207,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n206,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n205,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n204,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n203,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n202,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n201,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n200,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n199,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n198,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n197,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n196,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n195,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n194,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n193,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n192,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n191,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n190,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n290,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n289,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n288,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n287,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n286,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n285,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n284,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n283,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n282,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n281,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n280,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n279,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n278,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n277,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n276,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n275,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n274,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n273,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n272,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n271,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n270,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n269,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n268,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n267,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n266,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n265,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n264,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n263,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n262,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n261,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n260,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n259,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n258,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n257,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n256,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n255,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n254,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n253,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n252,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n251,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n250,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n249,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n248,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n247,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n246,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n245,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n244,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n243,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n242,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n241,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n240,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n239,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n238,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n237,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n236,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n235,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n234,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n233,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n232,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n231,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n230,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n229,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n228,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n227,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n226,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n225,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n224,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n286,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n285,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n284,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n283,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n282,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n281,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n280,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n279,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n278,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n277,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n276,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n275,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n274,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n273,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n272,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n271,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n270,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n269,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n268,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n267,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n266,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n265,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n264,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n263,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n262,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n261,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n260,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n259,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n258,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n257,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n256,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n255,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n254,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n253,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n252,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n251,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n250,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n249,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n248,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n247,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n246,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n245,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n244,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n243,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n242,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n241,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n240,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n239,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n238,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n237,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n236,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n235,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n234,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n233,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n232,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n231,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n230,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n229,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n228,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n227,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n226,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n225,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n224,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n223,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n222,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n221,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n220,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n219,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n218,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n217,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n283,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n282,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n281,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n280,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n279,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n278,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n277,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n276,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n275,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n274,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n273,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n272,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n271,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n270,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n269,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n268,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n267,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n266,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n265,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n264,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n263,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n262,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n261,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n260,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n259,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n258,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n257,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n256,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n255,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n254,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n253,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n252,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n251,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n250,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n249,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n248,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n247,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n246,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n245,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n244,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n243,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n242,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n241,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n240,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n239,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n238,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n237,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n236,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n235,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n234,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n233,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n232,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n231,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n230,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n229,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n228,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n227,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n226,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n225,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n224,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n223,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n222,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n221,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n220,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n219,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n218,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n217,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n216,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n215,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n283,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n282,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n281,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n280,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n279,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n278,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n277,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n276,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n275,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n274,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n273,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n272,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n271,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n270,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n269,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n268,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n267,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n266,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n265,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n264,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n263,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n262,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n261,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n260,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n259,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n258,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n257,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n256,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n255,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n254,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n253,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n252,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n251,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n250,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n249,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n248,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n247,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n246,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n245,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n244,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n243,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n242,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n241,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n240,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n239,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n238,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n237,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n236,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n235,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n234,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n233,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n232,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n231,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n230,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n229,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n228,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n227,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n226,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n225,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n224,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n223,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n222,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n280,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n279,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n278,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n277,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n276,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n275,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n274,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n273,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n272,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n271,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n270,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n269,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n268,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n267,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n266,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n265,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n264,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n263,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n262,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n261,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n260,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n259,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n258,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n257,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n256,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n255,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n254,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n253,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n252,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n251,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n250,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n249,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n248,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n247,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n246,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n245,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n244,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n243,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n242,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n241,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n240,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n239,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n238,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n237,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n236,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n235,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n234,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n233,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n232,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n231,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n230,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n229,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n228,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n227,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n226,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n225,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n224,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n223,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n222,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n221,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n220,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n219,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n218,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n217,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n216,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n215,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n279,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n278,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n277,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n276,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n275,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n274,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n273,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n272,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n271,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n270,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n269,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n268,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n267,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n266,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n265,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n264,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n263,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n262,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n261,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n260,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n259,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n258,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n257,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n256,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n255,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n254,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n253,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n252,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n251,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n250,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n249,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n248,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n247,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n246,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n245,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n244,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n243,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n242,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n241,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n240,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n239,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n238,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n237,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n236,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n235,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n234,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n233,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n232,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n231,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n230,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n229,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n228,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n227,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n226,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n225,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n224,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n223,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n222,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n221,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n220,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n219,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n218,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n217,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n216,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n215,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n214,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n240,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n239,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n238,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n237,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n236,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n235,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n234,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n233,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n232,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n231,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n230,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n229,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n228,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n227,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n226,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n225,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n224,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n223,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n222,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n221,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n220,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n219,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n218,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n217,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n216,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n215,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n214,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n213,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n212,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n211,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n210,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n209,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n208,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n207,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n206,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n205,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n204,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n203,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n202,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n201,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n200,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n199,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n198,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n197,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n196,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n195,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n194,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n193,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n192,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n191,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n190,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n290,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n289,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n288,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n287,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n286,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n285,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n284,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n283,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n282,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n281,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n280,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n279,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n278,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n277,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n276,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n275,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n274,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n273,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n272,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n271,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n270,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n269,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n268,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n267,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n266,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n265,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n264,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n263,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n262,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n261,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n260,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n259,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n258,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n257,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n256,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n255,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n254,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n253,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n252,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n251,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n250,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n249,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n248,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n247,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n246,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n245,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n244,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n243,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n242,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n241,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n240,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n239,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n238,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n237,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n236,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n235,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n234,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n233,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n232,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n231,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n230,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n229,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n228,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n227,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n226,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n225,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n224,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n286,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n285,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n284,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n283,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n282,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n281,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n280,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n279,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n278,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n277,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n276,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n275,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n274,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n273,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n272,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n271,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n270,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n269,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n268,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n267,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n266,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n265,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n264,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n263,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n262,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n261,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n260,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n259,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n258,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n257,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n256,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n255,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n254,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n253,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n252,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n251,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n250,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n249,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n248,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n247,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n246,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n245,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n244,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n243,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n242,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n241,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n240,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n239,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n238,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n237,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n236,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n235,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n234,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n233,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n232,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n231,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n230,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n229,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n228,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n227,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n226,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n225,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n224,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n223,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n222,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n221,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n220,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n219,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n218,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n217,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n283,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n282,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n281,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n280,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n279,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n278,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n277,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n276,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n275,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n274,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n273,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n272,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n271,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n270,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n269,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n268,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n267,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n266,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n265,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n264,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n263,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n262,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n261,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n260,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n259,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n258,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n257,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n256,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n255,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n254,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n253,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n252,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n251,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n250,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n249,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n248,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n247,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n246,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n245,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n244,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n243,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n242,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n241,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n240,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n239,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n238,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n237,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n236,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n235,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n234,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n233,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n232,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n231,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n230,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n229,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n228,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n227,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n226,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n225,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n224,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n223,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n222,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n221,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n220,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n219,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n218,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n217,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n216,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n215,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n283,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n282,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n281,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n280,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n279,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n278,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n277,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n276,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n275,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n274,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n273,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n272,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n271,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n270,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n269,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n268,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n267,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n266,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n265,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n264,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n263,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n262,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n261,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n260,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n259,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n258,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n257,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n256,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n255,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n254,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n253,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n252,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n251,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n250,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n249,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n248,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n247,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n246,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n245,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n244,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n243,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n242,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n241,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n240,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n239,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n238,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n237,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n236,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n235,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n234,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n233,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n232,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n231,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n230,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n229,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n228,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n227,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n226,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n225,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n224,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n223,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n222,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n280,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n279,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n278,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n277,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n276,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n275,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n274,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n273,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n272,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n271,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n270,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n269,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n268,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n267,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n266,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n265,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n264,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n263,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n262,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n261,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n260,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n259,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n258,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n257,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n256,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n255,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n254,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n253,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n252,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n251,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n250,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n249,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n248,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n247,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n246,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n245,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n244,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n243,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n242,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n241,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n240,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n239,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n238,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n237,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n236,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n235,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n234,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n233,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n232,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n231,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n230,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n229,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n228,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n227,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n226,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n225,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n224,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n223,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n222,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n221,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n220,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n219,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n218,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n217,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n216,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n215,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n279,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n278,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n277,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n276,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n275,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n274,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n273,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n272,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n271,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n270,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n269,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n268,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n267,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n266,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n265,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n264,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n263,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n262,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n261,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n260,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n259,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n258,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n257,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n256,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n255,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n254,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n253,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n252,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n251,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n250,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n249,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n248,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n247,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n246,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n245,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n244,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n243,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n242,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n241,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n240,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n239,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n238,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n237,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n236,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n235,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n234,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n233,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n232,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n231,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n230,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n229,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n228,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n227,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n226,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n225,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n224,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n223,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n222,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n221,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n220,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n219,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n218,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n217,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n216,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n215,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n214,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n240,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n239,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n238,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n237,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n236,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n235,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n234,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n233,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n232,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n231,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n230,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n229,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n228,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n227,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n226,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n225,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n224,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n223,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n222,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n221,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n220,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n219,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n218,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n217,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n216,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n215,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n214,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n213,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n212,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n211,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n210,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n209,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n208,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n207,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n206,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n205,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n204,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n203,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n202,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n201,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n200,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n199,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n198,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n197,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n196,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n195,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n194,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n193,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n192,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n191,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n190,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n290,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n289,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n288,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n287,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n286,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n285,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n284,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n283,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n282,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n281,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n280,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n279,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n278,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n277,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n276,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n275,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n274,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n273,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n272,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n271,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n270,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n269,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n268,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n267,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n266,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n265,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n264,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n263,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n262,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n261,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n260,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n259,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n258,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n257,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n256,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n255,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n254,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n253,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n252,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n251,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n250,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n249,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n248,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n247,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n246,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n245,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n244,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n243,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n242,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n241,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n240,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n239,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n238,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n237,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n236,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n235,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n234,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n233,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n232,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n231,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n230,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n229,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n228,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n227,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n226,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n225,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n224,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n286,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n285,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n284,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n283,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n282,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n281,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n280,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n279,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n278,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n277,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n276,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n275,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n274,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n273,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n272,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n271,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n270,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n269,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n268,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n267,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n266,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n265,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n264,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n263,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n262,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n261,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n260,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n259,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n258,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n257,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n256,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n255,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n254,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n253,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n252,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n251,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n250,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n249,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n248,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n247,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n246,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n245,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n244,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n243,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n242,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n241,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n240,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n239,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n238,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n237,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n236,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n235,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n234,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n233,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n232,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n231,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n230,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n229,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n228,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n227,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n226,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n225,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n224,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n223,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n222,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n221,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n220,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n219,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n218,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n217,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n283,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n282,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n281,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n280,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n279,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n278,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n277,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n276,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n275,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n274,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n273,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n272,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n271,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n270,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n269,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n268,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n267,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n266,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n265,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n264,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n263,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n262,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n261,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n260,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n259,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n258,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n257,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n256,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n255,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n254,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n253,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n252,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n251,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n250,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n249,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n248,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n247,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n246,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n245,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n244,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n243,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n242,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n241,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n240,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n239,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n238,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n237,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n236,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n235,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n234,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n233,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n232,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n231,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n230,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n229,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n228,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n227,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n226,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n225,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n224,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n223,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n222,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n221,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n220,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n219,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n218,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n217,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n216,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n215,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n283,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n282,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n281,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n280,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n279,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n278,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n277,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n276,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n275,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n274,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n273,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n272,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n271,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n270,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n269,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n268,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n267,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n266,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n265,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n264,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n263,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n262,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n261,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n260,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n259,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n258,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n257,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n256,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n255,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n254,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n253,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n252,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n251,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n250,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n249,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n248,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n247,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n246,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n245,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n244,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n243,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n242,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n241,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n240,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n239,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n238,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n237,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n236,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n235,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n234,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n233,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n232,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n231,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n230,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n229,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n228,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n227,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n226,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n225,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n224,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n223,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n222,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n280,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n279,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n278,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n277,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n276,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n275,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n274,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n273,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n272,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n271,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n270,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n269,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n268,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n267,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n266,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n265,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n264,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n263,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n262,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n261,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n260,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n259,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n258,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n257,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n256,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n255,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n254,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n253,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n252,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n251,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n250,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n249,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n248,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n247,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n246,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n245,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n244,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n243,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n242,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n241,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n240,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n239,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n238,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n237,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n236,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n235,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n234,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n233,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n232,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n231,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n230,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n229,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n228,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n227,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n226,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n225,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n224,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n223,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n222,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n221,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n220,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n219,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n218,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n217,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n216,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n215,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n279,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n278,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n277,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n276,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n275,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n274,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n273,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n272,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n271,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n270,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n269,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n268,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n267,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n266,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n265,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n264,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n263,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n262,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n261,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n260,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n259,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n258,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n257,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n256,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n255,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n254,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n253,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n252,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n251,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n250,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n249,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n248,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n247,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n246,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n245,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n244,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n243,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n242,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n241,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n240,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n239,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n238,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n237,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n236,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n235,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n234,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n233,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n232,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n231,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n230,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n229,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n228,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n227,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n226,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n225,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n224,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n223,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n222,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n221,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n220,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n219,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n218,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n217,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n216,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n215,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n214,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n240,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n239,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n238,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n237,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n236,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n235,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n234,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n233,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n232,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n231,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n230,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n229,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n228,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n227,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n226,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n225,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n224,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n223,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n222,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n221,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n220,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n219,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n218,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n217,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n216,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n215,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n214,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n213,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n212,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n211,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n210,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n209,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n208,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n207,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n206,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n205,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n204,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n203,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n202,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n201,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n200,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n199,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n198,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n197,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n196,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n195,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n194,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n193,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n192,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n191,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n190,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n290,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n289,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n288,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n287,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n286,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n285,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n284,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n283,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n282,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n281,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n280,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n279,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n278,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n277,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n276,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n275,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n274,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n273,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n272,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n271,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n270,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n269,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n268,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n267,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n266,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n265,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n264,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n263,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n262,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n261,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n260,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n259,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n258,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n257,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n256,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n255,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n254,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n253,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n252,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n251,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n250,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n249,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n248,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n247,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n246,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n245,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n244,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n243,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n242,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n241,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n240,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n239,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n238,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n237,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n236,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n235,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n234,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n233,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n232,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n231,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n230,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n229,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n228,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n227,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n226,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n225,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n224,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n286,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n285,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n284,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n283,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n282,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n281,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n280,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n279,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n278,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n277,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n276,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n275,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n274,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n273,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n272,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n271,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n270,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n269,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n268,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n267,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n266,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n265,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n264,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n263,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n262,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n261,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n260,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n259,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n258,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n257,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n256,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n255,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n254,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n253,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n252,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n251,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n250,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n249,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n248,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n247,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n246,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n245,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n244,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n243,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n242,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n241,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n240,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n239,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n238,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n237,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n236,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n235,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n234,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n233,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n232,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n231,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n230,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n229,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n228,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n227,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n226,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n225,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n224,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n223,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n222,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n221,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n220,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n219,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n218,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n217,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n283,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n282,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n281,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n280,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n279,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n278,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n277,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n276,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n275,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n274,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n273,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n272,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n271,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n270,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n269,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n268,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n267,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n266,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n265,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n264,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n263,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n262,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n261,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n260,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n259,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n258,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n257,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n256,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n255,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n254,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n253,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n252,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n251,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n250,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n249,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n248,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n247,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n246,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n245,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n244,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n243,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n242,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n241,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n240,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n239,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n238,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n237,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n236,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n235,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n234,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n233,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n232,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n231,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n230,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n229,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n228,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n227,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n226,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n225,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n224,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n223,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n222,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n221,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n220,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n219,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n218,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n217,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n216,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n215,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n283,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n282,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n281,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n280,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n279,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n278,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n277,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n276,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n275,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n274,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n273,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n272,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n271,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n270,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n269,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n268,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n267,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n266,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n265,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n264,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n263,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n262,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n261,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n260,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n259,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n258,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n257,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n256,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n255,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n254,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n253,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n252,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n251,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n250,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n249,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n248,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n247,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n246,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n245,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n244,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n243,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n242,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n241,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n240,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n239,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n238,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n237,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n236,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n235,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n234,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n233,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n232,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n231,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n230,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n229,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n228,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n227,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n226,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n225,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n224,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n223,
         F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n222,
         K0K1_KeyMUX_And_Red_KeyMUX_n89, K0K1_KeyMUX_And_Red_KeyMUX_n88,
         K0K1_KeyMUX_And_Red_KeyMUX_n87, K0K1_KeyMUX_And_Red_KeyMUX_n86,
         K0K1_KeyMUX_And_Red_KeyMUX_n85, K0K1_KeyMUX_And_Red_KeyMUX_n84,
         K0K1_KeyMUX_And_Red_KeyMUX_n83, K0K1_KeyMUX_And_Red_KeyMUX_n82,
         K0K1_KeyMUX_And_Red_KeyMUX_n81, K0K1_KeyMUX_And_Red_KeyMUX_n80,
         K0K1_KeyMUX_And_Red_KeyMUX_n79, K0K1_KeyMUX_And_Red_KeyMUX_n78,
         K0K1_KeyMUX_And_Red_KeyMUX_n77, K0K1_KeyMUX_And_Red_KeyMUX_n76,
         K0K1_KeyMUX_And_Red_KeyMUX_n75, K0K1_KeyMUX_And_Red_KeyMUX_n74,
         K0K1_KeyMUX_And_Red_KeyMUX_n73, K0K1_KeyMUX_And_Red_KeyMUX_n72,
         K0K1_KeyMUX_And_Red_KeyMUX_n71, K0K1_KeyMUX_And_Red_KeyMUX_n70,
         K0K1_KeyMUX_And_Red_KeyMUX_n69, K0K1_KeyMUX_And_Red_KeyMUX_n68,
         K0K1_KeyMUX_And_Red_KeyMUX_n67, K0K1_KeyMUX_And_Red_KeyMUX_n66,
         K0K1_KeyMUX_And_Red_KeyMUX_n65, K0K1_KeyMUX_And_Red_KeyMUX_n64,
         K0K1_KeyMUX_And_Red_KeyMUX_n63, K0K1_KeyMUX_And_Red_KeyMUX_n62,
         K0K1_KeyMUX_And_Red_KeyMUX_n61, K0K1_KeyMUX_And_Red_KeyMUX_n60,
         K0K1_KeyMUX_And_Red_KeyMUX_n59, K0K1_KeyMUX_And_Red_KeyMUX_n58,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_0_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_0_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_0_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_0_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_0_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_0_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_0_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_0_n23,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_1_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_1_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_1_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_1_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_1_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_1_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_1_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_1_n23,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_2_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_2_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_2_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_2_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_2_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_2_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_2_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_2_n23,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_3_n31,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_3_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_3_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_3_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_3_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_3_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_3_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_3_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_4_n31,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_4_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_4_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_4_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_4_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_4_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_4_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_4_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_5_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_5_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_5_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_5_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_5_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_5_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_5_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_5_n23,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_6_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_6_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_6_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_6_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_6_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_6_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_6_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_6_n23,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_7_n31,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_7_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_7_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_7_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_7_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_7_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_7_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_7_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_8_n31,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_8_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_8_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_8_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_8_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_8_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_8_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_8_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_9_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_9_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_9_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_9_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_9_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_9_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_9_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_9_n23,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_10_n31,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_10_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_10_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_10_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_10_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_10_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_10_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_10_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_11_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_11_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_11_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_11_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_11_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_11_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_11_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_11_n23,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_12_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_12_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_12_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_12_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_12_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_12_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_12_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_12_n23,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_13_n31,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_13_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_13_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_13_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_13_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_13_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_13_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_13_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_14_n31,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_14_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_14_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_14_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_14_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_14_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_14_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_14_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_15_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_15_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_15_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_15_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_15_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_15_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_15_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_15_n23,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_16_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_16_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_16_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_16_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_16_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_16_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_16_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_16_n23,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_17_n31,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_17_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_17_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_17_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_17_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_17_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_17_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_17_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_18_n31,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_18_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_18_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_18_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_18_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_18_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_18_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_18_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_19_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_19_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_19_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_19_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_19_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_19_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_19_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_19_n23,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_20_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_20_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_20_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_20_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_20_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_20_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_20_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_20_n23,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_21_n31,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_21_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_21_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_21_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_21_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_21_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_21_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_21_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_22_n31,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_22_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_22_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_22_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_22_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_22_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_22_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_22_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_23_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_23_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_23_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_23_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_23_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_23_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_23_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_23_n23,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_24_n31,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_24_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_24_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_24_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_24_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_24_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_24_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_24_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_25_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_25_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_25_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_25_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_25_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_25_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_25_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_25_n23,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_26_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_26_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_26_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_26_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_26_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_26_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_26_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_26_n23,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_27_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_27_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_27_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_27_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_27_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_27_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_27_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_27_n23,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_28_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_28_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_28_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_28_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_28_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_28_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_28_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_28_n23,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_29_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_29_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_29_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_29_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_29_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_29_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_29_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_29_n23,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_30_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_30_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_30_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_30_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_30_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_30_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_30_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_30_n23,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_31_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_31_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_31_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_31_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_31_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_31_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_31_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_31_n23,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_32_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_32_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_32_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_32_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_32_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_32_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_32_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_32_n23,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_33_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_33_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_33_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_33_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_33_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_33_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_33_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_33_n23,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_34_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_34_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_34_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_34_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_34_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_34_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_34_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_34_n23,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_35_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_35_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_35_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_35_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_35_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_35_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_35_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_35_n23,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_36_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_36_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_36_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_36_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_36_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_36_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_36_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_36_n23,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_37_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_37_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_37_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_37_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_37_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_37_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_37_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_37_n23,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_38_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_38_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_38_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_38_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_38_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_38_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_38_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_38_n23,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_39_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_39_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_39_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_39_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_39_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_39_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_39_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_39_n23,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_40_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_40_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_40_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_40_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_40_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_40_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_40_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_40_n23,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_41_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_41_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_41_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_41_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_41_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_41_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_41_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_41_n23,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_42_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_42_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_42_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_42_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_42_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_42_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_42_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_42_n23,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_43_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_43_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_43_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_43_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_43_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_43_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_43_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_43_n23,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_44_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_44_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_44_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_44_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_44_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_44_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_44_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_44_n23,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_45_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_45_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_45_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_45_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_45_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_45_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_45_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_45_n23,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_46_n31,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_46_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_46_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_46_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_46_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_46_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_46_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_46_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_47_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_47_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_47_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_47_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_47_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_47_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_47_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_47_n23,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_48_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_48_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_48_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_48_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_48_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_48_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_48_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_48_n23,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_49_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_49_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_49_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_49_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_49_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_49_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_49_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_49_n23,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_50_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_50_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_50_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_50_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_50_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_50_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_50_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_50_n23,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_51_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_51_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_51_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_51_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_51_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_51_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_51_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_51_n23,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_52_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_52_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_52_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_52_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_52_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_52_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_52_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_52_n23,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_53_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_53_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_53_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_53_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_53_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_53_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_53_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_53_n23,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_54_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_54_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_54_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_54_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_54_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_54_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_54_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_54_n23,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_55_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_55_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_55_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_55_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_55_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_55_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_55_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_55_n23,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_56_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_56_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_56_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_56_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_56_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_56_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_56_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_56_n23,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_57_n31,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_57_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_57_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_57_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_57_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_57_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_57_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_57_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_58_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_58_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_58_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_58_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_58_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_58_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_58_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_58_n23,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_59_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_59_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_59_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_59_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_59_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_59_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_59_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_59_n23,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_60_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_60_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_60_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_60_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_60_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_60_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_60_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_60_n23,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_61_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_61_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_61_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_61_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_61_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_61_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_61_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_61_n23,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_62_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_62_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_62_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_62_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_62_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_62_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_62_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_62_n23,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_63_n31,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_63_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_63_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_63_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_63_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_63_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_63_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_63_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_64_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_64_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_64_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_64_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_64_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_64_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_64_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_64_n23,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_65_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_65_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_65_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_65_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_65_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_65_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_65_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_65_n23,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_66_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_66_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_66_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_66_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_66_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_66_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_66_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_66_n23,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_67_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_67_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_67_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_67_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_67_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_67_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_67_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_67_n23,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_68_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_68_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_68_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_68_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_68_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_68_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_68_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_68_n23,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_69_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_69_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_69_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_69_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_69_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_69_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_69_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_69_n23,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_70_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_70_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_70_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_70_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_70_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_70_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_70_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_70_n23,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_71_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_71_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_71_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_71_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_71_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_71_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_71_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_71_n23,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_72_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_72_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_72_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_72_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_72_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_72_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_72_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_72_n23,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_73_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_73_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_73_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_73_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_73_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_73_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_73_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_73_n23,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_74_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_74_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_74_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_74_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_74_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_74_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_74_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_74_n23,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_75_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_75_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_75_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_75_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_75_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_75_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_75_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_75_n23,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_76_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_76_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_76_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_76_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_76_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_76_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_76_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_76_n23,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_77_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_77_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_77_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_77_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_77_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_77_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_77_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_77_n23,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_78_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_78_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_78_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_78_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_78_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_78_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_78_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_78_n23,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_79_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_79_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_79_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_79_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_79_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_79_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_79_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_79_n23,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_80_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_80_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_80_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_80_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_80_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_80_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_80_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_80_n23,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_81_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_81_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_81_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_81_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_81_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_81_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_81_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_81_n23,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_82_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_82_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_82_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_82_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_82_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_82_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_82_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_82_n23,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_83_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_83_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_83_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_83_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_83_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_83_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_83_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_83_n23,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_84_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_84_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_84_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_84_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_84_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_84_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_84_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_84_n23,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_85_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_85_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_85_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_85_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_85_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_85_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_85_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_85_n23,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_86_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_86_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_86_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_86_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_86_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_86_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_86_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_86_n23,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_87_n31,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_87_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_87_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_87_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_87_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_87_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_87_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_87_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_88_n31,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_88_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_88_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_88_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_88_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_88_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_88_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_88_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_89_n31,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_89_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_89_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_89_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_89_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_89_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_89_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_89_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_90_n31,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_90_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_90_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_90_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_90_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_90_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_90_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_90_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_91_n31,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_91_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_91_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_91_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_91_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_91_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_91_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_91_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_92_n31,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_92_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_92_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_92_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_92_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_92_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_92_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_92_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_93_n31,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_93_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_93_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_93_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_93_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_93_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_93_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_93_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_94_n31,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_94_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_94_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_94_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_94_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_94_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_94_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_94_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_95_n32,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_95_n31,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_95_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_95_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_95_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_95_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_95_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_95_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_96_n32,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_96_n31,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_96_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_96_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_96_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_96_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_96_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_96_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_97_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_97_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_97_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_97_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_97_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_97_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_97_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_97_n23,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_98_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_98_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_98_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_98_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_98_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_98_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_98_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_98_n23,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_99_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_99_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_99_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_99_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_99_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_99_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_99_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_99_n23,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_100_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_100_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_100_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_100_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_100_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_100_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_100_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_100_n23,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_101_n31,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_101_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_101_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_101_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_101_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_101_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_101_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_101_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_102_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_102_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_102_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_102_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_102_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_102_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_102_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_102_n23,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_103_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_103_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_103_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_103_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_103_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_103_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_103_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_103_n23,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_104_n31,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_104_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_104_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_104_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_104_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_104_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_104_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_104_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_105_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_105_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_105_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_105_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_105_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_105_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_105_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_105_n23,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_106_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_106_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_106_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_106_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_106_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_106_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_106_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_106_n23,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_107_n31,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_107_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_107_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_107_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_107_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_107_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_107_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_107_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_108_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_108_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_108_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_108_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_108_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_108_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_108_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_108_n23,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_109_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_109_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_109_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_109_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_109_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_109_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_109_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_109_n23,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_110_n31,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_110_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_110_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_110_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_110_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_110_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_110_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_110_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_111_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_111_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_111_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_111_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_111_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_111_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_111_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_111_n23,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_112_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_112_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_112_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_112_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_112_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_112_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_112_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_112_n23,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_113_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_113_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_113_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_113_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_113_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_113_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_113_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_113_n23,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_114_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_114_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_114_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_114_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_114_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_114_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_114_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_114_n23,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_115_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_115_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_115_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_115_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_115_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_115_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_115_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_115_n23,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_116_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_116_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_116_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_116_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_116_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_116_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_116_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_116_n23,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_117_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_117_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_117_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_117_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_117_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_117_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_117_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_117_n23,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_118_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_118_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_118_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_118_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_118_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_118_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_118_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_118_n23,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_119_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_119_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_119_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_119_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_119_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_119_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_119_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_119_n23,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_120_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_120_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_120_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_120_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_120_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_120_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_120_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_120_n23,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_121_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_121_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_121_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_121_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_121_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_121_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_121_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_121_n23,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_122_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_122_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_122_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_122_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_122_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_122_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_122_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_122_n23,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_123_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_123_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_123_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_123_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_123_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_123_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_123_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_123_n23,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_124_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_124_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_124_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_124_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_124_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_124_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_124_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_124_n23,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_125_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_125_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_125_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_125_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_125_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_125_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_125_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_125_n23,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_126_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_126_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_126_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_126_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_126_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_126_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_126_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_126_n23,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_127_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_127_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_127_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_127_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_127_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_127_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_127_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_127_n23,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_128_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_128_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_128_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_128_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_128_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_128_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_128_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_128_n23,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_129_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_129_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_129_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_129_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_129_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_129_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_129_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_129_n23,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_130_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_130_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_130_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_130_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_130_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_130_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_130_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_130_n23,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_131_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_131_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_131_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_131_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_131_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_131_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_131_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_131_n23,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_132_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_132_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_132_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_132_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_132_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_132_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_132_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_132_n23,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_133_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_133_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_133_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_133_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_133_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_133_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_133_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_133_n23,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_134_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_134_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_134_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_134_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_134_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_134_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_134_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_134_n23,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_135_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_135_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_135_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_135_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_135_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_135_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_135_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_135_n23,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_136_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_136_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_136_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_136_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_136_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_136_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_136_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_136_n23,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_137_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_137_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_137_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_137_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_137_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_137_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_137_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_137_n23,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_138_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_138_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_138_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_138_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_138_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_138_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_138_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_138_n23,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_139_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_139_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_139_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_139_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_139_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_139_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_139_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_139_n23,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_140_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_140_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_140_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_140_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_140_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_140_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_140_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_140_n23,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_141_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_141_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_141_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_141_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_141_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_141_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_141_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_141_n23,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_142_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_142_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_142_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_142_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_142_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_142_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_142_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_142_n23,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_143_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_143_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_143_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_143_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_143_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_143_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_143_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_143_n23,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_144_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_144_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_144_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_144_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_144_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_144_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_144_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_144_n23,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_145_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_145_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_145_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_145_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_145_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_145_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_145_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_145_n23,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_146_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_146_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_146_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_146_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_146_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_146_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_146_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_146_n23,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_147_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_147_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_147_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_147_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_147_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_147_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_147_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_147_n23,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_148_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_148_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_148_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_148_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_148_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_148_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_148_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_148_n23,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_149_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_149_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_149_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_149_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_149_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_149_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_149_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_149_n23,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_150_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_150_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_150_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_150_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_150_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_150_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_150_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_150_n23,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_151_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_151_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_151_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_151_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_151_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_151_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_151_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_151_n23,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_152_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_152_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_152_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_152_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_152_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_152_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_152_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_152_n23,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_153_n31,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_153_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_153_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_153_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_153_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_153_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_153_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_153_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_154_n31,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_154_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_154_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_154_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_154_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_154_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_154_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_154_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_155_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_155_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_155_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_155_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_155_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_155_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_155_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_155_n23,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_156_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_156_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_156_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_156_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_156_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_156_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_156_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_156_n23,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_157_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_157_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_157_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_157_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_157_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_157_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_157_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_157_n23,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_158_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_158_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_158_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_158_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_158_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_158_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_158_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_158_n23,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_159_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_159_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_159_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_159_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_159_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_159_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_159_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_159_n23,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_160_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_160_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_160_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_160_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_160_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_160_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_160_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_160_n23,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_161_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_161_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_161_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_161_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_161_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_161_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_161_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_161_n23,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_162_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_162_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_162_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_162_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_162_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_162_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_162_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_162_n23,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_163_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_163_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_163_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_163_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_163_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_163_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_163_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_163_n23,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_164_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_164_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_164_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_164_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_164_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_164_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_164_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_164_n23,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_165_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_165_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_165_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_165_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_165_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_165_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_165_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_165_n23,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_166_n31,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_166_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_166_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_166_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_166_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_166_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_166_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_166_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_167_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_167_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_167_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_167_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_167_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_167_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_167_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_167_n23,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_168_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_168_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_168_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_168_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_168_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_168_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_168_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_168_n23,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_169_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_169_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_169_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_169_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_169_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_169_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_169_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_169_n23,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_170_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_170_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_170_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_170_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_170_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_170_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_170_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_170_n23,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_171_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_171_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_171_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_171_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_171_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_171_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_171_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_171_n23,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_172_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_172_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_172_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_172_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_172_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_172_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_172_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_172_n23,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_173_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_173_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_173_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_173_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_173_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_173_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_173_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_173_n23,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_174_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_174_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_174_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_174_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_174_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_174_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_174_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_174_n23,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_175_n30,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_175_n29,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_175_n28,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_175_n27,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_175_n26,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_175_n25,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_175_n24,
         K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_175_n23,
         Red_K0Inst_LFInst_0_LFInst_0_n3, Red_K0Inst_LFInst_0_LFInst_1_n3,
         Red_K0Inst_LFInst_1_LFInst_0_n3, Red_K0Inst_LFInst_1_LFInst_1_n3,
         Red_K0Inst_LFInst_2_LFInst_0_n3, Red_K0Inst_LFInst_2_LFInst_1_n3,
         Red_K0Inst_LFInst_3_LFInst_0_n3, Red_K0Inst_LFInst_3_LFInst_1_n3,
         Red_K0Inst_LFInst_4_LFInst_0_n3, Red_K0Inst_LFInst_4_LFInst_1_n3,
         Red_K0Inst_LFInst_5_LFInst_0_n3, Red_K0Inst_LFInst_5_LFInst_1_n3,
         Red_K0Inst_LFInst_6_LFInst_0_n3, Red_K0Inst_LFInst_6_LFInst_1_n3,
         Red_K0Inst_LFInst_7_LFInst_0_n3, Red_K0Inst_LFInst_7_LFInst_1_n3,
         Red_K0Inst_LFInst_8_LFInst_0_n3, Red_K0Inst_LFInst_8_LFInst_1_n3,
         Red_K0Inst_LFInst_9_LFInst_0_n3, Red_K0Inst_LFInst_9_LFInst_1_n3,
         Red_K0Inst_LFInst_10_LFInst_0_n3, Red_K0Inst_LFInst_10_LFInst_1_n3,
         Red_K0Inst_LFInst_11_LFInst_0_n3, Red_K0Inst_LFInst_11_LFInst_1_n3,
         Red_K0Inst_LFInst_12_LFInst_0_n3, Red_K0Inst_LFInst_12_LFInst_1_n3,
         Red_K0Inst_LFInst_13_LFInst_0_n3, Red_K0Inst_LFInst_13_LFInst_1_n3,
         Red_K0Inst_LFInst_14_LFInst_0_n3, Red_K0Inst_LFInst_14_LFInst_1_n3,
         Red_K0Inst_LFInst_15_LFInst_0_n3, Red_K0Inst_LFInst_15_LFInst_1_n3,
         Red_K1Inst_LFInst_0_LFInst_0_n3, Red_K1Inst_LFInst_0_LFInst_1_n3,
         Red_K1Inst_LFInst_1_LFInst_0_n3, Red_K1Inst_LFInst_1_LFInst_1_n3,
         Red_K1Inst_LFInst_2_LFInst_0_n3, Red_K1Inst_LFInst_2_LFInst_1_n3,
         Red_K1Inst_LFInst_3_LFInst_0_n3, Red_K1Inst_LFInst_3_LFInst_1_n3,
         Red_K1Inst_LFInst_4_LFInst_0_n3, Red_K1Inst_LFInst_4_LFInst_1_n3,
         Red_K1Inst_LFInst_5_LFInst_0_n3, Red_K1Inst_LFInst_5_LFInst_1_n3,
         Red_K1Inst_LFInst_6_LFInst_0_n3, Red_K1Inst_LFInst_6_LFInst_1_n3,
         Red_K1Inst_LFInst_7_LFInst_0_n3, Red_K1Inst_LFInst_7_LFInst_1_n3,
         Red_K1Inst_LFInst_8_LFInst_0_n3, Red_K1Inst_LFInst_8_LFInst_1_n3,
         Red_K1Inst_LFInst_9_LFInst_0_n3, Red_K1Inst_LFInst_9_LFInst_1_n3,
         Red_K1Inst_LFInst_10_LFInst_0_n3, Red_K1Inst_LFInst_10_LFInst_1_n3,
         Red_K1Inst_LFInst_11_LFInst_0_n3, Red_K1Inst_LFInst_11_LFInst_1_n3,
         Red_K1Inst_LFInst_12_LFInst_0_n3, Red_K1Inst_LFInst_12_LFInst_1_n3,
         Red_K1Inst_LFInst_13_LFInst_0_n3, Red_K1Inst_LFInst_13_LFInst_1_n3,
         Red_K1Inst_LFInst_14_LFInst_0_n3, Red_K1Inst_LFInst_14_LFInst_1_n3,
         Red_K1Inst_LFInst_15_LFInst_0_n3, Red_K1Inst_LFInst_15_LFInst_1_n3,
         FSMMUX_MUXInst_1_n4, FSMMUX_MUXInst_2_n4, FSMMUX_MUXInst_4_n4,
         FSMMUX_MUXInst_5_n4, FSMMUX_MUXInst_6_n4,
         F_FSM_Inst_LFInst_0_LFInst_0_n3, F_FSM_Inst_LFInst_1_LFInst_0_n3,
         F_FSM_Inst_LFInst_1_LFInst_1_n3, F_SD1_StateUpdate_Done_Inst_n5,
         F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_0_n12,
         F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_0_n11,
         F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_0_n10,
         F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_0_n9,
         F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_0_n8,
         F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_0_n6,
         F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_0_n5,
         F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_0_n4,
         F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_1_n13,
         F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_1_n12,
         F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_1_n11,
         F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_1_n10,
         F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_1_n9,
         F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_1_n8,
         F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_1_n7,
         F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_1_n6,
         F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_1_n5,
         F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_1_n4,
         F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_1_n3,
         F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_1_n2,
         F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_1_n1,
         F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_2_n15,
         F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_2_n14,
         F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_2_n13,
         F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_2_n12,
         F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_2_n11,
         F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_2_n10,
         F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_2_n9,
         F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_2_n8,
         F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_2_n7,
         F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_2_n6,
         F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_2_n5,
         F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_2_n3,
         F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_2_n2,
         F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_2_n1,
         F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_inst_3_n14,
         F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_inst_3_n13,
         F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_inst_3_n12,
         F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_inst_3_n11,
         F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_inst_3_n10,
         F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_inst_3_n9,
         F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_inst_3_n8,
         F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_inst_3_n7,
         F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_inst_3_n6,
         F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_inst_3_n5,
         F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_inst_3_n4,
         F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_inst_4_n12,
         F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_inst_4_n11,
         F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_inst_4_n10,
         F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_inst_4_n9,
         F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_inst_4_n7,
         F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_inst_4_n6,
         F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_inst_4_n5,
         F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_inst_4_n4,
         F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_inst_4_n3,
         F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_inst_4_n2,
         F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_inst_4_n1,
         F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_inst_5_n12,
         F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_inst_5_n11,
         F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_inst_5_n10,
         F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_inst_5_n9,
         F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_inst_5_n8,
         F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_inst_5_n7,
         F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_inst_5_n6,
         F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_inst_5_n5,
         F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_inst_5_n4,
         F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_inst_5_n3,
         F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_inst_5_n2,
         F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_inst_5_n1,
         F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_6_n17,
         F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_6_n16,
         F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_6_n15,
         F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_6_n14,
         F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_6_n13,
         F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_6_n12,
         F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_6_n11,
         F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_6_n10,
         F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_6_n9,
         F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_6_n8,
         F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_6_n7,
         F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_6_n6,
         F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_6_n5,
         F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_6_n4,
         F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_6_n3,
         F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_6_n2,
         F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_6_n1,
         F_SD1_SelectsUpdate_Bit0_Inst_n11, F_SD1_SelectsUpdate_Bit0_Inst_n10,
         F_SD1_SelectsUpdate_Bit0_Inst_n9, F_SD1_SelectsUpdate_Bit0_Inst_n8,
         F_SD1_SelectsUpdate_Bit0_Inst_n7, F_SD1_SelectsUpdate_Bit0_Inst_n6,
         F_SD1_SelectsUpdate_Bit0_Inst_n5, F_SD1_SelectsUpdate_Bit0_Inst_n4,
         F_SD1_SelectsUpdate_Bit0_Inst_n3, Red_FSMMUX_MUXInst_4_n4,
         Red_FSMMUX_MUXInst_5_n4, Red_FSMMUX_MUXInst_6_n4,
         Red_FSMMUX_MUXInst_11_n4, Red_FSMMUX_MUXInst_12_n4,
         Red_FSMMUX_MUXInst_13_n4, F_SD2_RedStateUpdate_Done_Inst_n9,
         F_SD2_RedStateUpdate_Done_Inst_n8, F_SD2_RedStateUpdate_Done_Inst_n7,
         F_SD2_RedStateUpdate_Done_Inst_n6, F_SD2_RedStateUpdate_Done_Inst_n5,
         F_SD2_RedStateUpdate_Done_Inst_n4, F_SD2_RedStateUpdate_Done_Inst_n3,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n329,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n328,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n327,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n326,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n325,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n324,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n323,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n322,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n321,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n320,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n319,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n318,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n317,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n316,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n315,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n314,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n313,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n312,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n311,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n310,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n309,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n308,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n307,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n306,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n305,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n304,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n303,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n302,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n301,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n300,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n299,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n298,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n297,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n296,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n295,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n294,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n293,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n292,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n291,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n290,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n289,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n288,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n287,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n286,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n285,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n284,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n283,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n282,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n281,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n280,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n279,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n278,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n277,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n276,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n275,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n274,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n273,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n272,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n271,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n270,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n269,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n268,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n267,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n266,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n265,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n264,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n263,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n262,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n261,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n260,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n259,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n258,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n257,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n256,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n255,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n254,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n253,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n252,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n251,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n250,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n249,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n248,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n247,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n246,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n245,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n244,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n243,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n242,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n241,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n240,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n239,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n238,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n237,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n236,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n235,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n234,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n233,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n232,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n231,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n230,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n229,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n228,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n227,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n226,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n225,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n224,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n223,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n222,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n221,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n220,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n219,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n218,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n217,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n216,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n215,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n214,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n213,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n212,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n211,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n210,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n209,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n208,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n207,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n206,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n205,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n204,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n203,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n202,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n201,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n200,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n199,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n198,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n197,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n196,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n195,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n317,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n316,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n315,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n314,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n313,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n312,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n311,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n310,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n309,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n308,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n307,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n306,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n305,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n304,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n303,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n302,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n301,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n300,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n299,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n298,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n297,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n296,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n295,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n294,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n293,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n292,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n291,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n290,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n289,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n288,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n287,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n286,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n285,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n284,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n283,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n282,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n281,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n280,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n279,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n278,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n277,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n276,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n275,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n274,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n273,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n272,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n271,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n270,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n269,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n268,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n267,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n266,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n265,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n264,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n263,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n262,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n261,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n260,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n259,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n258,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n257,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n256,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n255,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n254,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n253,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n252,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n251,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n250,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n249,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n248,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n247,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n246,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n245,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n244,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n243,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n242,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n241,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n240,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n239,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n238,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n237,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n236,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n235,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n234,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n233,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n232,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n231,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n230,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n229,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n228,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n227,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n226,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n225,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n224,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n223,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n222,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n221,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n220,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n219,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n218,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n217,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n216,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n215,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n214,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n213,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n212,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n211,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n210,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n209,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n208,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n207,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n206,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n205,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n204,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n203,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n202,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n201,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n200,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n199,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n198,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n197,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n196,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n195,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n194,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_n233,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_n232,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_n231,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_n230,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_n229,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_n228,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_n227,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_n226,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_n225,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_n224,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_n223,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_n222,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_n221,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_n220,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_n219,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_n218,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_n217,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_n216,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_n215,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_n214,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_n213,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_n212,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_n211,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_n210,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_n209,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_n208,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_n207,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_n206,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_n205,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_n204,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_n203,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_n202,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_n201,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_n200,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_n199,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_n198,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_n197,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_n196,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_n195,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_n228,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_n227,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_n226,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_n225,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_n224,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_n223,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_n222,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_n221,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_n220,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_n219,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_n218,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_n217,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_n216,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_n215,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_n214,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_n213,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_n212,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_n211,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_n210,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_n209,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_n208,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_n207,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_n206,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_n205,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_n204,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_n203,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_n202,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_n201,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_n200,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_n199,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_n198,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_n197,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_n196,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_n195,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_n194,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_4_n71,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_4_n70,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_4_n69,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_4_n68,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_4_n67,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_4_n66,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_4_n65,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_4_n64,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_4_n63,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_4_n62,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_4_n61,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_4_n60,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_4_n59,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_4_n58,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_4_n57,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_4_n56,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_4_n55,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_4_n54,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_4_n53,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_4_n52,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_4_n51,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_4_n50,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_4_n49,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_4_n48,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_4_n47,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n125,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n124,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n123,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n122,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n121,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n120,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n119,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n118,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n117,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n116,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n115,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n114,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n113,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n112,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n111,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n110,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n109,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n108,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n107,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n106,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n105,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n104,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n103,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n102,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n101,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n100,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n99,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n98,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n97,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n96,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n95,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n94,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n93,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n92,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n91,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n90,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n89,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n88,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n87,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n86,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n85,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n84,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n83,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n82,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n81,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n80,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n79,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n78,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n77,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n76,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n75,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n74,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n73,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n151,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n150,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n149,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n148,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n147,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n146,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n145,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n144,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n143,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n142,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n141,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n140,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n139,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n138,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n137,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n136,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n135,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n134,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n133,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n132,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n131,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n130,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n129,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n128,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n127,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n126,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n125,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n124,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n123,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n122,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n121,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n120,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n119,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n118,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n117,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n116,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n115,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n114,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n113,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n112,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n111,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n110,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n109,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n108,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n107,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n106,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n105,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n104,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n103,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n102,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n101,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n100,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n99,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n98,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n97,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n96,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n95,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n94,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n93,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n92,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n91,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n90,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n89,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n88,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n87,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n140,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n139,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n138,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n137,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n136,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n135,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n134,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n133,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n132,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n131,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n130,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n129,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n128,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n127,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n126,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n125,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n124,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n123,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n122,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n121,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n120,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n119,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n118,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n117,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n116,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n115,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n114,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n113,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n112,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n111,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n110,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n109,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n108,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n107,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n106,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n105,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n104,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n103,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n102,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n101,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n100,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n99,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n98,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n97,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n96,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n95,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_8_n108,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_8_n107,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_8_n106,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_8_n105,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_8_n104,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_8_n103,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_8_n102,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_8_n101,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_8_n100,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_8_n99,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_8_n98,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_8_n97,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_8_n96,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_8_n95,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_8_n94,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_8_n93,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_8_n92,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_8_n91,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_8_n90,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_8_n89,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_8_n88,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_8_n87,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_8_n86,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_8_n85,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_8_n84,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_8_n83,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_9_n119,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_9_n118,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_9_n117,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_9_n116,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_9_n115,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_9_n114,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_9_n113,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_9_n112,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_9_n111,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_9_n110,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_9_n109,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_9_n108,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_9_n107,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_9_n106,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_9_n105,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_9_n104,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_9_n103,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_9_n102,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_9_n101,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_9_n100,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_9_n99,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_9_n98,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_9_n97,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_9_n96,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_9_n95,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_9_n94,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_9_n93,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_9_n92,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_9_n91,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_9_n90,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n130,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n129,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n128,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n127,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n126,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n125,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n124,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n123,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n122,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n121,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n120,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n119,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n118,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n117,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n116,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n115,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n114,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n113,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n112,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n111,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n110,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n109,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n108,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n107,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n106,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n105,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n104,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n103,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n102,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n101,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n100,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n99,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n98,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n97,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n96,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n95,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n94,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n93,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n92,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n91,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n90,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n89,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n88,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n87,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n124,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n123,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n122,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n121,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n120,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n119,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n118,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n117,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n116,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n115,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n114,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n113,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n112,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n111,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n110,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n109,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n108,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n107,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n106,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n105,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n104,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n103,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n102,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n101,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n100,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n99,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n98,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n97,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n96,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n95,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n94,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n93,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n92,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n91,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n90,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n89,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n88,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n87,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n86,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n85,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n84,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n83,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_12_n111,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_12_n110,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_12_n109,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_12_n108,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_12_n107,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_12_n106,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_12_n105,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_12_n104,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_12_n103,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_12_n102,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_12_n101,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_12_n100,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_12_n99,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_12_n98,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_12_n97,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_12_n96,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_12_n95,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_12_n94,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_12_n93,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_12_n92,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_12_n91,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_12_n90,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_12_n89,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_12_n88,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_12_n87,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_12_n86,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_12_n85,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_12_n84,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_13_n96,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_13_n95,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_13_n94,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_13_n93,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_13_n92,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_13_n91,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_13_n90,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_13_n89,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_13_n88,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_13_n87,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_13_n86,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_13_n85,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_13_n84,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_13_n83,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_13_n82,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_13_n81,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_13_n80,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_13_n79,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_13_n78,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_13_n77,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_13_n76,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_13_n75,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_13_n74,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_13_n73,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_13_n72,
         F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_13_n71,
         Red_selectsMUX_MUXInst_0_n4, Red_selectsMUX_MUXInst_1_n4,
         Red_selectsMUX_MUXInst_2_n6, Red_selectsMUX_MUXInst_2_n5,
         Red_selectsMUX_MUXInst_3_n4,
         F_SD2_Red_SelectsUpdate_Inst_F_SD2_Red_SelectsUpdate_Bit_Inst_0_n12,
         F_SD2_Red_SelectsUpdate_Inst_F_SD2_Red_SelectsUpdate_Bit_Inst_0_n11,
         F_SD2_Red_SelectsUpdate_Inst_F_SD2_Red_SelectsUpdate_Bit_Inst_0_n10,
         F_SD2_Red_SelectsUpdate_Inst_F_SD2_Red_SelectsUpdate_Bit_Inst_0_n9,
         F_SD2_Red_SelectsUpdate_Inst_F_SD2_Red_SelectsUpdate_Bit_Inst_0_n8,
         F_SD2_Red_SelectsUpdate_Inst_F_SD2_Red_SelectsUpdate_Bit_Inst_0_n7,
         F_SD2_Red_SelectsUpdate_Inst_F_SD2_Red_SelectsUpdate_Bit_Inst_0_n6,
         F_SD2_Red_SelectsUpdate_Inst_F_SD2_Red_SelectsUpdate_Bit_Inst_1_n12,
         F_SD2_Red_SelectsUpdate_Inst_F_SD2_Red_SelectsUpdate_Bit_Inst_1_n11,
         F_SD2_Red_SelectsUpdate_Inst_F_SD2_Red_SelectsUpdate_Bit_Inst_1_n10,
         F_SD2_Red_SelectsUpdate_Inst_F_SD2_Red_SelectsUpdate_Bit_Inst_1_n9,
         F_SD2_Red_SelectsUpdate_Inst_F_SD2_Red_SelectsUpdate_Bit_Inst_1_n8,
         F_SD2_Red_SelectsUpdate_Inst_F_SD2_Red_SelectsUpdate_Bit_Inst_1_n7,
         F_SD2_Red_SelectsUpdate_Inst_F_SD2_Red_SelectsUpdate_Bit_Inst_1_n6,
         F_SD2_Red_SelectsUpdate_Inst_F_SD2_Red_SelectsUpdate_Bit_Inst_2_n29,
         F_SD2_Red_SelectsUpdate_Inst_F_SD2_Red_SelectsUpdate_Bit_Inst_2_n28,
         F_SD2_Red_SelectsUpdate_Inst_F_SD2_Red_SelectsUpdate_Bit_Inst_2_n27,
         F_SD2_Red_SelectsUpdate_Inst_F_SD2_Red_SelectsUpdate_Bit_Inst_2_n26,
         F_SD2_Red_SelectsUpdate_Inst_F_SD2_Red_SelectsUpdate_Bit_Inst_2_n25,
         F_SD2_Red_SelectsUpdate_Inst_F_SD2_Red_SelectsUpdate_Bit_Inst_2_n24,
         F_SD2_Red_SelectsUpdate_Inst_F_SD2_Red_SelectsUpdate_Bit_Inst_2_n23,
         F_SD2_Red_SelectsUpdate_Inst_F_SD2_Red_SelectsUpdate_Bit_Inst_3_n12,
         F_SD2_Red_SelectsUpdate_Inst_F_SD2_Red_SelectsUpdate_Bit_Inst_3_n11,
         F_SD2_Red_SelectsUpdate_Inst_F_SD2_Red_SelectsUpdate_Bit_Inst_3_n10,
         F_SD2_Red_SelectsUpdate_Inst_F_SD2_Red_SelectsUpdate_Bit_Inst_3_n9,
         F_SD2_Red_SelectsUpdate_Inst_F_SD2_Red_SelectsUpdate_Bit_Inst_3_n8,
         F_SD2_Red_SelectsUpdate_Inst_F_SD2_Red_SelectsUpdate_Bit_Inst_3_n7,
         F_SD2_Red_SelectsUpdate_Inst_F_SD2_Red_SelectsUpdate_Bit_Inst_3_n6,
         Output_MUX_n10, Output_MUX_n9, Output_MUX_n8, Output_MUX_n7;
  wire   [63:0] Feedback;
  wire   [63:32] MCInput;
  wire   [63:0] MCOutput;
  wire   [63:0] AddRoundKeyOutput;
  wire   [7:0] RoundConstant;
  wire   [63:0] StateRegOutput;
  wire   [111:0] StateRegOutputF;
  wire   [111:0] Red_StateRegOutput;
  wire   [111:0] CipherErrorVec;
  wire   [63:0] OutputRegIn;
  wire   [111:0] Red_Input;
  wire   [111:0] Red_Feedback;
  wire   [111:56] Red_MCInput;
  wire   [111:0] Red_MCOutput;
  wire   [111:0] Red_AddRoundKeyOutput;
  wire   [13:0] Red_RoundConstant;
  wire   [4:0] KeyMux_sel_input;
  wire   [111:0] KeyMux_D0_input;
  wire   [111:0] KeyMux_D1_input;
  wire   [63:0] SelectedKey;
  wire   [111:0] Red_SelectedKey;
  wire   [6:0] FSMReg;
  wire   [6:3] FSM;
  wire   [13:0] FSMF;
  wire   [13:0] FSMErrorVec;
  wire   [6:2] FSMUpdate;
  wire   [13:0] Red_FSMReg;
  wire   [1:0] Red_done;
  wire   [13:0] Red_FSMUpdate;
  wire   [3:0] Red_selectsReg;
  wire   [3:0] Red_selectsNext;

  BUF_X2 U3 ( .A(KeyMux_sel_input[1]), .Z(n6) );
  BUF_X1 U4 ( .A(KeyMux_sel_input[4]), .Z(n7) );
  BUF_X1 U5 ( .A(KeyMux_sel_input[0]), .Z(n5) );
  MUX2_X1 InputMUX_MUXInst_0_U1 ( .A(Feedback[0]), .B(Input[0]), .S(rst), .Z(
        MCOutput[0]) );
  MUX2_X1 InputMUX_MUXInst_1_U1 ( .A(Feedback[1]), .B(Input[1]), .S(rst), .Z(
        MCOutput[1]) );
  MUX2_X1 InputMUX_MUXInst_2_U1 ( .A(Feedback[2]), .B(Input[2]), .S(rst), .Z(
        MCOutput[2]) );
  MUX2_X1 InputMUX_MUXInst_3_U1 ( .A(Feedback[3]), .B(Input[3]), .S(rst), .Z(
        MCOutput[3]) );
  MUX2_X1 InputMUX_MUXInst_4_U1 ( .A(Feedback[4]), .B(Input[4]), .S(rst), .Z(
        MCOutput[4]) );
  MUX2_X1 InputMUX_MUXInst_5_U1 ( .A(Feedback[5]), .B(Input[5]), .S(rst), .Z(
        MCOutput[5]) );
  MUX2_X1 InputMUX_MUXInst_6_U1 ( .A(Feedback[6]), .B(Input[6]), .S(rst), .Z(
        MCOutput[6]) );
  MUX2_X1 InputMUX_MUXInst_7_U1 ( .A(Feedback[7]), .B(Input[7]), .S(rst), .Z(
        MCOutput[7]) );
  MUX2_X1 InputMUX_MUXInst_8_U1 ( .A(Feedback[8]), .B(Input[8]), .S(rst), .Z(
        MCOutput[8]) );
  MUX2_X1 InputMUX_MUXInst_9_U1 ( .A(Feedback[9]), .B(Input[9]), .S(rst), .Z(
        MCOutput[9]) );
  MUX2_X1 InputMUX_MUXInst_10_U1 ( .A(Feedback[10]), .B(Input[10]), .S(rst), 
        .Z(MCOutput[10]) );
  MUX2_X1 InputMUX_MUXInst_11_U1 ( .A(Feedback[11]), .B(Input[11]), .S(rst), 
        .Z(MCOutput[11]) );
  MUX2_X1 InputMUX_MUXInst_12_U1 ( .A(Feedback[12]), .B(Input[12]), .S(rst), 
        .Z(MCOutput[12]) );
  MUX2_X1 InputMUX_MUXInst_13_U1 ( .A(Feedback[13]), .B(Input[13]), .S(rst), 
        .Z(MCOutput[13]) );
  MUX2_X1 InputMUX_MUXInst_14_U1 ( .A(Feedback[14]), .B(Input[14]), .S(rst), 
        .Z(MCOutput[14]) );
  MUX2_X1 InputMUX_MUXInst_15_U1 ( .A(Feedback[15]), .B(Input[15]), .S(rst), 
        .Z(MCOutput[15]) );
  MUX2_X1 InputMUX_MUXInst_16_U1 ( .A(Feedback[16]), .B(Input[16]), .S(rst), 
        .Z(MCOutput[16]) );
  MUX2_X1 InputMUX_MUXInst_17_U1 ( .A(Feedback[17]), .B(Input[17]), .S(rst), 
        .Z(MCOutput[17]) );
  MUX2_X1 InputMUX_MUXInst_18_U1 ( .A(Feedback[18]), .B(Input[18]), .S(rst), 
        .Z(MCOutput[18]) );
  MUX2_X1 InputMUX_MUXInst_19_U1 ( .A(Feedback[19]), .B(Input[19]), .S(rst), 
        .Z(MCOutput[19]) );
  MUX2_X1 InputMUX_MUXInst_20_U1 ( .A(Feedback[20]), .B(Input[20]), .S(rst), 
        .Z(MCOutput[20]) );
  MUX2_X1 InputMUX_MUXInst_21_U1 ( .A(Feedback[21]), .B(Input[21]), .S(rst), 
        .Z(MCOutput[21]) );
  MUX2_X1 InputMUX_MUXInst_22_U1 ( .A(Feedback[22]), .B(Input[22]), .S(rst), 
        .Z(MCOutput[22]) );
  MUX2_X1 InputMUX_MUXInst_23_U1 ( .A(Feedback[23]), .B(Input[23]), .S(rst), 
        .Z(MCOutput[23]) );
  MUX2_X1 InputMUX_MUXInst_24_U1 ( .A(Feedback[24]), .B(Input[24]), .S(rst), 
        .Z(MCOutput[24]) );
  MUX2_X1 InputMUX_MUXInst_25_U1 ( .A(Feedback[25]), .B(Input[25]), .S(rst), 
        .Z(MCOutput[25]) );
  MUX2_X1 InputMUX_MUXInst_26_U1 ( .A(Feedback[26]), .B(Input[26]), .S(rst), 
        .Z(MCOutput[26]) );
  MUX2_X1 InputMUX_MUXInst_27_U1 ( .A(Feedback[27]), .B(Input[27]), .S(rst), 
        .Z(MCOutput[27]) );
  MUX2_X1 InputMUX_MUXInst_28_U1 ( .A(Feedback[28]), .B(Input[28]), .S(rst), 
        .Z(MCOutput[28]) );
  MUX2_X1 InputMUX_MUXInst_29_U1 ( .A(Feedback[29]), .B(Input[29]), .S(rst), 
        .Z(MCOutput[29]) );
  MUX2_X1 InputMUX_MUXInst_30_U1 ( .A(Feedback[30]), .B(Input[30]), .S(rst), 
        .Z(MCOutput[30]) );
  MUX2_X1 InputMUX_MUXInst_31_U1 ( .A(Feedback[31]), .B(Input[31]), .S(rst), 
        .Z(MCOutput[31]) );
  MUX2_X1 InputMUX_MUXInst_32_U1 ( .A(Feedback[32]), .B(Input[32]), .S(rst), 
        .Z(MCInput[32]) );
  MUX2_X1 InputMUX_MUXInst_33_U1 ( .A(Feedback[33]), .B(Input[33]), .S(rst), 
        .Z(MCInput[33]) );
  MUX2_X1 InputMUX_MUXInst_34_U1 ( .A(Feedback[34]), .B(Input[34]), .S(rst), 
        .Z(MCInput[34]) );
  MUX2_X1 InputMUX_MUXInst_35_U1 ( .A(Feedback[35]), .B(Input[35]), .S(rst), 
        .Z(MCInput[35]) );
  MUX2_X1 InputMUX_MUXInst_36_U1 ( .A(Feedback[36]), .B(Input[36]), .S(rst), 
        .Z(MCInput[36]) );
  MUX2_X1 InputMUX_MUXInst_37_U1 ( .A(Feedback[37]), .B(Input[37]), .S(rst), 
        .Z(MCInput[37]) );
  MUX2_X1 InputMUX_MUXInst_38_U1 ( .A(Feedback[38]), .B(Input[38]), .S(rst), 
        .Z(MCInput[38]) );
  MUX2_X1 InputMUX_MUXInst_39_U1 ( .A(Feedback[39]), .B(Input[39]), .S(rst), 
        .Z(MCInput[39]) );
  MUX2_X1 InputMUX_MUXInst_40_U1 ( .A(Feedback[40]), .B(Input[40]), .S(rst), 
        .Z(MCInput[40]) );
  MUX2_X1 InputMUX_MUXInst_41_U1 ( .A(Feedback[41]), .B(Input[41]), .S(rst), 
        .Z(MCInput[41]) );
  MUX2_X1 InputMUX_MUXInst_42_U1 ( .A(Feedback[42]), .B(Input[42]), .S(rst), 
        .Z(MCInput[42]) );
  MUX2_X1 InputMUX_MUXInst_43_U1 ( .A(Feedback[43]), .B(Input[43]), .S(rst), 
        .Z(MCInput[43]) );
  MUX2_X1 InputMUX_MUXInst_44_U1 ( .A(Feedback[44]), .B(Input[44]), .S(rst), 
        .Z(MCInput[44]) );
  MUX2_X1 InputMUX_MUXInst_45_U1 ( .A(Feedback[45]), .B(Input[45]), .S(rst), 
        .Z(MCInput[45]) );
  MUX2_X1 InputMUX_MUXInst_46_U1 ( .A(Feedback[46]), .B(Input[46]), .S(rst), 
        .Z(MCInput[46]) );
  MUX2_X1 InputMUX_MUXInst_47_U1 ( .A(Feedback[47]), .B(Input[47]), .S(rst), 
        .Z(MCInput[47]) );
  MUX2_X1 InputMUX_MUXInst_48_U1 ( .A(Feedback[48]), .B(Input[48]), .S(rst), 
        .Z(MCInput[48]) );
  MUX2_X1 InputMUX_MUXInst_49_U1 ( .A(Feedback[49]), .B(Input[49]), .S(rst), 
        .Z(MCInput[49]) );
  MUX2_X1 InputMUX_MUXInst_50_U1 ( .A(Feedback[50]), .B(Input[50]), .S(rst), 
        .Z(MCInput[50]) );
  MUX2_X1 InputMUX_MUXInst_51_U1 ( .A(Feedback[51]), .B(Input[51]), .S(rst), 
        .Z(MCInput[51]) );
  MUX2_X1 InputMUX_MUXInst_52_U1 ( .A(Feedback[52]), .B(Input[52]), .S(rst), 
        .Z(MCInput[52]) );
  MUX2_X1 InputMUX_MUXInst_53_U1 ( .A(Feedback[53]), .B(Input[53]), .S(rst), 
        .Z(MCInput[53]) );
  MUX2_X1 InputMUX_MUXInst_54_U1 ( .A(Feedback[54]), .B(Input[54]), .S(rst), 
        .Z(MCInput[54]) );
  MUX2_X1 InputMUX_MUXInst_55_U1 ( .A(Feedback[55]), .B(Input[55]), .S(rst), 
        .Z(MCInput[55]) );
  MUX2_X1 InputMUX_MUXInst_56_U1 ( .A(Feedback[56]), .B(Input[56]), .S(rst), 
        .Z(MCInput[56]) );
  MUX2_X1 InputMUX_MUXInst_57_U1 ( .A(Feedback[57]), .B(Input[57]), .S(rst), 
        .Z(MCInput[57]) );
  MUX2_X1 InputMUX_MUXInst_58_U1 ( .A(Feedback[58]), .B(Input[58]), .S(rst), 
        .Z(MCInput[58]) );
  MUX2_X1 InputMUX_MUXInst_59_U1 ( .A(Feedback[59]), .B(Input[59]), .S(rst), 
        .Z(MCInput[59]) );
  MUX2_X1 InputMUX_MUXInst_60_U1 ( .A(Feedback[60]), .B(Input[60]), .S(rst), 
        .Z(MCInput[60]) );
  MUX2_X1 InputMUX_MUXInst_61_U1 ( .A(Feedback[61]), .B(Input[61]), .S(rst), 
        .Z(MCInput[61]) );
  MUX2_X1 InputMUX_MUXInst_62_U1 ( .A(Feedback[62]), .B(Input[62]), .S(rst), 
        .Z(MCInput[62]) );
  MUX2_X1 InputMUX_MUXInst_63_U1 ( .A(Feedback[63]), .B(Input[63]), .S(rst), 
        .Z(MCInput[63]) );
  XNOR2_X1 MCInst_XOR_r0_Inst_0_U2 ( .A(MCInst_XOR_r0_Inst_0_n5), .B(
        MCOutput[16]), .ZN(MCOutput[48]) );
  XNOR2_X1 MCInst_XOR_r0_Inst_0_U1 ( .A(MCOutput[0]), .B(MCInput[48]), .ZN(
        MCInst_XOR_r0_Inst_0_n5) );
  XOR2_X1 MCInst_XOR_r1_Inst_0_U1 ( .A(MCInput[32]), .B(MCOutput[0]), .Z(
        MCOutput[32]) );
  XNOR2_X1 MCInst_XOR_r0_Inst_1_U2 ( .A(MCInst_XOR_r0_Inst_1_n5), .B(
        MCOutput[17]), .ZN(MCOutput[49]) );
  XNOR2_X1 MCInst_XOR_r0_Inst_1_U1 ( .A(MCOutput[1]), .B(MCInput[49]), .ZN(
        MCInst_XOR_r0_Inst_1_n5) );
  XOR2_X1 MCInst_XOR_r1_Inst_1_U1 ( .A(MCInput[33]), .B(MCOutput[1]), .Z(
        MCOutput[33]) );
  XNOR2_X1 MCInst_XOR_r0_Inst_2_U2 ( .A(MCInst_XOR_r0_Inst_2_n5), .B(
        MCOutput[18]), .ZN(MCOutput[50]) );
  XNOR2_X1 MCInst_XOR_r0_Inst_2_U1 ( .A(MCOutput[2]), .B(MCInput[50]), .ZN(
        MCInst_XOR_r0_Inst_2_n5) );
  XOR2_X1 MCInst_XOR_r1_Inst_2_U1 ( .A(MCInput[34]), .B(MCOutput[2]), .Z(
        MCOutput[34]) );
  XNOR2_X1 MCInst_XOR_r0_Inst_3_U2 ( .A(MCInst_XOR_r0_Inst_3_n5), .B(
        MCOutput[19]), .ZN(MCOutput[51]) );
  XNOR2_X1 MCInst_XOR_r0_Inst_3_U1 ( .A(MCOutput[3]), .B(MCInput[51]), .ZN(
        MCInst_XOR_r0_Inst_3_n5) );
  XOR2_X1 MCInst_XOR_r1_Inst_3_U1 ( .A(MCInput[35]), .B(MCOutput[3]), .Z(
        MCOutput[35]) );
  XNOR2_X1 MCInst_XOR_r0_Inst_4_U2 ( .A(MCInst_XOR_r0_Inst_4_n5), .B(
        MCOutput[20]), .ZN(MCOutput[52]) );
  XNOR2_X1 MCInst_XOR_r0_Inst_4_U1 ( .A(MCOutput[4]), .B(MCInput[52]), .ZN(
        MCInst_XOR_r0_Inst_4_n5) );
  XOR2_X1 MCInst_XOR_r1_Inst_4_U1 ( .A(MCInput[36]), .B(MCOutput[4]), .Z(
        MCOutput[36]) );
  XNOR2_X1 MCInst_XOR_r0_Inst_5_U2 ( .A(MCInst_XOR_r0_Inst_5_n5), .B(
        MCOutput[21]), .ZN(MCOutput[53]) );
  XNOR2_X1 MCInst_XOR_r0_Inst_5_U1 ( .A(MCOutput[5]), .B(MCInput[53]), .ZN(
        MCInst_XOR_r0_Inst_5_n5) );
  XOR2_X1 MCInst_XOR_r1_Inst_5_U1 ( .A(MCInput[37]), .B(MCOutput[5]), .Z(
        MCOutput[37]) );
  XNOR2_X1 MCInst_XOR_r0_Inst_6_U2 ( .A(MCInst_XOR_r0_Inst_6_n5), .B(
        MCOutput[22]), .ZN(MCOutput[54]) );
  XNOR2_X1 MCInst_XOR_r0_Inst_6_U1 ( .A(MCOutput[6]), .B(MCInput[54]), .ZN(
        MCInst_XOR_r0_Inst_6_n5) );
  XOR2_X1 MCInst_XOR_r1_Inst_6_U1 ( .A(MCInput[38]), .B(MCOutput[6]), .Z(
        MCOutput[38]) );
  XNOR2_X1 MCInst_XOR_r0_Inst_7_U2 ( .A(MCInst_XOR_r0_Inst_7_n5), .B(
        MCOutput[23]), .ZN(MCOutput[55]) );
  XNOR2_X1 MCInst_XOR_r0_Inst_7_U1 ( .A(MCOutput[7]), .B(MCInput[55]), .ZN(
        MCInst_XOR_r0_Inst_7_n5) );
  XOR2_X1 MCInst_XOR_r1_Inst_7_U1 ( .A(MCInput[39]), .B(MCOutput[7]), .Z(
        MCOutput[39]) );
  XNOR2_X1 MCInst_XOR_r0_Inst_8_U2 ( .A(MCInst_XOR_r0_Inst_8_n5), .B(
        MCOutput[24]), .ZN(MCOutput[56]) );
  XNOR2_X1 MCInst_XOR_r0_Inst_8_U1 ( .A(MCOutput[8]), .B(MCInput[56]), .ZN(
        MCInst_XOR_r0_Inst_8_n5) );
  XOR2_X1 MCInst_XOR_r1_Inst_8_U1 ( .A(MCInput[40]), .B(MCOutput[8]), .Z(
        MCOutput[40]) );
  XNOR2_X1 MCInst_XOR_r0_Inst_9_U2 ( .A(MCInst_XOR_r0_Inst_9_n5), .B(
        MCOutput[25]), .ZN(MCOutput[57]) );
  XNOR2_X1 MCInst_XOR_r0_Inst_9_U1 ( .A(MCOutput[9]), .B(MCInput[57]), .ZN(
        MCInst_XOR_r0_Inst_9_n5) );
  XOR2_X1 MCInst_XOR_r1_Inst_9_U1 ( .A(MCInput[41]), .B(MCOutput[9]), .Z(
        MCOutput[41]) );
  XNOR2_X1 MCInst_XOR_r0_Inst_10_U2 ( .A(MCInst_XOR_r0_Inst_10_n5), .B(
        MCOutput[26]), .ZN(MCOutput[58]) );
  XNOR2_X1 MCInst_XOR_r0_Inst_10_U1 ( .A(MCOutput[10]), .B(MCInput[58]), .ZN(
        MCInst_XOR_r0_Inst_10_n5) );
  XOR2_X1 MCInst_XOR_r1_Inst_10_U1 ( .A(MCInput[42]), .B(MCOutput[10]), .Z(
        MCOutput[42]) );
  XNOR2_X1 MCInst_XOR_r0_Inst_11_U2 ( .A(MCInst_XOR_r0_Inst_11_n5), .B(
        MCOutput[27]), .ZN(MCOutput[59]) );
  XNOR2_X1 MCInst_XOR_r0_Inst_11_U1 ( .A(MCOutput[11]), .B(MCInput[59]), .ZN(
        MCInst_XOR_r0_Inst_11_n5) );
  XOR2_X1 MCInst_XOR_r1_Inst_11_U1 ( .A(MCInput[43]), .B(MCOutput[11]), .Z(
        MCOutput[43]) );
  XNOR2_X1 MCInst_XOR_r0_Inst_12_U2 ( .A(MCInst_XOR_r0_Inst_12_n5), .B(
        MCOutput[28]), .ZN(MCOutput[60]) );
  XNOR2_X1 MCInst_XOR_r0_Inst_12_U1 ( .A(MCOutput[12]), .B(MCInput[60]), .ZN(
        MCInst_XOR_r0_Inst_12_n5) );
  XOR2_X1 MCInst_XOR_r1_Inst_12_U1 ( .A(MCInput[44]), .B(MCOutput[12]), .Z(
        MCOutput[44]) );
  XNOR2_X1 MCInst_XOR_r0_Inst_13_U2 ( .A(MCInst_XOR_r0_Inst_13_n5), .B(
        MCOutput[29]), .ZN(MCOutput[61]) );
  XNOR2_X1 MCInst_XOR_r0_Inst_13_U1 ( .A(MCOutput[13]), .B(MCInput[61]), .ZN(
        MCInst_XOR_r0_Inst_13_n5) );
  XOR2_X1 MCInst_XOR_r1_Inst_13_U1 ( .A(MCInput[45]), .B(MCOutput[13]), .Z(
        MCOutput[45]) );
  XNOR2_X1 MCInst_XOR_r0_Inst_14_U2 ( .A(MCInst_XOR_r0_Inst_14_n5), .B(
        MCOutput[30]), .ZN(MCOutput[62]) );
  XNOR2_X1 MCInst_XOR_r0_Inst_14_U1 ( .A(MCOutput[14]), .B(MCInput[62]), .ZN(
        MCInst_XOR_r0_Inst_14_n5) );
  XOR2_X1 MCInst_XOR_r1_Inst_14_U1 ( .A(MCInput[46]), .B(MCOutput[14]), .Z(
        MCOutput[46]) );
  XNOR2_X1 MCInst_XOR_r0_Inst_15_U2 ( .A(MCInst_XOR_r0_Inst_15_n5), .B(
        MCOutput[31]), .ZN(MCOutput[63]) );
  XNOR2_X1 MCInst_XOR_r0_Inst_15_U1 ( .A(MCOutput[15]), .B(MCInput[63]), .ZN(
        MCInst_XOR_r0_Inst_15_n5) );
  XOR2_X1 MCInst_XOR_r1_Inst_15_U1 ( .A(MCInput[47]), .B(MCOutput[15]), .Z(
        MCOutput[47]) );
  XOR2_X1 AddKeyXOR1_XORInst_0_0_U1 ( .A(MCOutput[48]), .B(SelectedKey[48]), 
        .Z(AddRoundKeyOutput[48]) );
  XOR2_X1 AddKeyXOR1_XORInst_0_1_U1 ( .A(MCOutput[49]), .B(SelectedKey[49]), 
        .Z(AddRoundKeyOutput[49]) );
  XOR2_X1 AddKeyXOR1_XORInst_0_2_U1 ( .A(MCOutput[50]), .B(SelectedKey[50]), 
        .Z(AddRoundKeyOutput[50]) );
  XOR2_X1 AddKeyXOR1_XORInst_0_3_U1 ( .A(MCOutput[51]), .B(SelectedKey[51]), 
        .Z(AddRoundKeyOutput[51]) );
  XOR2_X1 AddKeyXOR1_XORInst_1_0_U1 ( .A(MCOutput[52]), .B(SelectedKey[52]), 
        .Z(AddRoundKeyOutput[52]) );
  XOR2_X1 AddKeyXOR1_XORInst_1_1_U1 ( .A(MCOutput[53]), .B(SelectedKey[53]), 
        .Z(AddRoundKeyOutput[53]) );
  XOR2_X1 AddKeyXOR1_XORInst_1_2_U1 ( .A(MCOutput[54]), .B(SelectedKey[54]), 
        .Z(AddRoundKeyOutput[54]) );
  XOR2_X1 AddKeyXOR1_XORInst_1_3_U1 ( .A(MCOutput[55]), .B(SelectedKey[55]), 
        .Z(AddRoundKeyOutput[55]) );
  XOR2_X1 AddKeyXOR1_XORInst_2_0_U1 ( .A(MCOutput[56]), .B(SelectedKey[56]), 
        .Z(AddRoundKeyOutput[56]) );
  XOR2_X1 AddKeyXOR1_XORInst_2_1_U1 ( .A(MCOutput[57]), .B(SelectedKey[57]), 
        .Z(AddRoundKeyOutput[57]) );
  XOR2_X1 AddKeyXOR1_XORInst_2_2_U1 ( .A(MCOutput[58]), .B(SelectedKey[58]), 
        .Z(AddRoundKeyOutput[58]) );
  XOR2_X1 AddKeyXOR1_XORInst_2_3_U1 ( .A(MCOutput[59]), .B(SelectedKey[59]), 
        .Z(AddRoundKeyOutput[59]) );
  XOR2_X1 AddKeyXOR1_XORInst_3_0_U1 ( .A(MCOutput[60]), .B(SelectedKey[60]), 
        .Z(AddRoundKeyOutput[60]) );
  XOR2_X1 AddKeyXOR1_XORInst_3_1_U1 ( .A(MCOutput[61]), .B(SelectedKey[61]), 
        .Z(AddRoundKeyOutput[61]) );
  XOR2_X1 AddKeyXOR1_XORInst_3_2_U1 ( .A(MCOutput[62]), .B(SelectedKey[62]), 
        .Z(AddRoundKeyOutput[62]) );
  XOR2_X1 AddKeyXOR1_XORInst_3_3_U1 ( .A(MCOutput[63]), .B(SelectedKey[63]), 
        .Z(AddRoundKeyOutput[63]) );
  XNOR2_X1 AddKeyConstXOR_XORInst_0_0_U2 ( .A(AddKeyConstXOR_XORInst_0_0_n5), 
        .B(SelectedKey[40]), .ZN(AddRoundKeyOutput[40]) );
  XNOR2_X1 AddKeyConstXOR_XORInst_0_0_U1 ( .A(RoundConstant[0]), .B(
        MCOutput[40]), .ZN(AddKeyConstXOR_XORInst_0_0_n5) );
  XNOR2_X1 AddKeyConstXOR_XORInst_0_1_U2 ( .A(AddKeyConstXOR_XORInst_0_1_n5), 
        .B(SelectedKey[41]), .ZN(AddRoundKeyOutput[41]) );
  XNOR2_X1 AddKeyConstXOR_XORInst_0_1_U1 ( .A(RoundConstant[1]), .B(
        MCOutput[41]), .ZN(AddKeyConstXOR_XORInst_0_1_n5) );
  XNOR2_X1 AddKeyConstXOR_XORInst_0_2_U2 ( .A(AddKeyConstXOR_XORInst_0_2_n5), 
        .B(SelectedKey[42]), .ZN(AddRoundKeyOutput[42]) );
  XNOR2_X1 AddKeyConstXOR_XORInst_0_2_U1 ( .A(RoundConstant[2]), .B(
        MCOutput[42]), .ZN(AddKeyConstXOR_XORInst_0_2_n5) );
  XOR2_X1 AddKeyConstXOR_XORInst_0_3_U1 ( .A(MCOutput[43]), .B(SelectedKey[43]), .Z(AddRoundKeyOutput[43]) );
  XNOR2_X1 AddKeyConstXOR_XORInst_1_0_U2 ( .A(AddKeyConstXOR_XORInst_1_0_n5), 
        .B(SelectedKey[44]), .ZN(AddRoundKeyOutput[44]) );
  XNOR2_X1 AddKeyConstXOR_XORInst_1_0_U1 ( .A(RoundConstant[4]), .B(
        MCOutput[44]), .ZN(AddKeyConstXOR_XORInst_1_0_n5) );
  XNOR2_X1 AddKeyConstXOR_XORInst_1_1_U2 ( .A(AddKeyConstXOR_XORInst_1_1_n5), 
        .B(SelectedKey[45]), .ZN(AddRoundKeyOutput[45]) );
  XNOR2_X1 AddKeyConstXOR_XORInst_1_1_U1 ( .A(RoundConstant[5]), .B(
        MCOutput[45]), .ZN(AddKeyConstXOR_XORInst_1_1_n5) );
  XNOR2_X1 AddKeyConstXOR_XORInst_1_2_U2 ( .A(AddKeyConstXOR_XORInst_1_2_n5), 
        .B(SelectedKey[46]), .ZN(AddRoundKeyOutput[46]) );
  XNOR2_X1 AddKeyConstXOR_XORInst_1_2_U1 ( .A(RoundConstant[6]), .B(
        MCOutput[46]), .ZN(AddKeyConstXOR_XORInst_1_2_n5) );
  XNOR2_X1 AddKeyConstXOR_XORInst_1_3_U2 ( .A(AddKeyConstXOR_XORInst_1_3_n5), 
        .B(SelectedKey[47]), .ZN(AddRoundKeyOutput[47]) );
  XNOR2_X1 AddKeyConstXOR_XORInst_1_3_U1 ( .A(RoundConstant[7]), .B(
        MCOutput[47]), .ZN(AddKeyConstXOR_XORInst_1_3_n5) );
  XOR2_X1 AddKeyXOR2_XORInst_0_0_U1 ( .A(MCOutput[0]), .B(SelectedKey[0]), .Z(
        AddRoundKeyOutput[0]) );
  XOR2_X1 AddKeyXOR2_XORInst_0_1_U1 ( .A(MCOutput[1]), .B(SelectedKey[1]), .Z(
        AddRoundKeyOutput[1]) );
  XOR2_X1 AddKeyXOR2_XORInst_0_2_U1 ( .A(MCOutput[2]), .B(SelectedKey[2]), .Z(
        AddRoundKeyOutput[2]) );
  XOR2_X1 AddKeyXOR2_XORInst_0_3_U1 ( .A(MCOutput[3]), .B(SelectedKey[3]), .Z(
        AddRoundKeyOutput[3]) );
  XOR2_X1 AddKeyXOR2_XORInst_1_0_U1 ( .A(MCOutput[4]), .B(SelectedKey[4]), .Z(
        AddRoundKeyOutput[4]) );
  XOR2_X1 AddKeyXOR2_XORInst_1_1_U1 ( .A(MCOutput[5]), .B(SelectedKey[5]), .Z(
        AddRoundKeyOutput[5]) );
  XOR2_X1 AddKeyXOR2_XORInst_1_2_U1 ( .A(MCOutput[6]), .B(SelectedKey[6]), .Z(
        AddRoundKeyOutput[6]) );
  XOR2_X1 AddKeyXOR2_XORInst_1_3_U1 ( .A(MCOutput[7]), .B(SelectedKey[7]), .Z(
        AddRoundKeyOutput[7]) );
  XOR2_X1 AddKeyXOR2_XORInst_2_0_U1 ( .A(MCOutput[8]), .B(SelectedKey[8]), .Z(
        AddRoundKeyOutput[8]) );
  XOR2_X1 AddKeyXOR2_XORInst_2_1_U1 ( .A(MCOutput[9]), .B(SelectedKey[9]), .Z(
        AddRoundKeyOutput[9]) );
  XOR2_X1 AddKeyXOR2_XORInst_2_2_U1 ( .A(MCOutput[10]), .B(SelectedKey[10]), 
        .Z(AddRoundKeyOutput[10]) );
  XOR2_X1 AddKeyXOR2_XORInst_2_3_U1 ( .A(MCOutput[11]), .B(SelectedKey[11]), 
        .Z(AddRoundKeyOutput[11]) );
  XOR2_X1 AddKeyXOR2_XORInst_3_0_U1 ( .A(MCOutput[12]), .B(SelectedKey[12]), 
        .Z(AddRoundKeyOutput[12]) );
  XOR2_X1 AddKeyXOR2_XORInst_3_1_U1 ( .A(MCOutput[13]), .B(SelectedKey[13]), 
        .Z(AddRoundKeyOutput[13]) );
  XOR2_X1 AddKeyXOR2_XORInst_3_2_U1 ( .A(MCOutput[14]), .B(SelectedKey[14]), 
        .Z(AddRoundKeyOutput[14]) );
  XOR2_X1 AddKeyXOR2_XORInst_3_3_U1 ( .A(MCOutput[15]), .B(SelectedKey[15]), 
        .Z(AddRoundKeyOutput[15]) );
  XOR2_X1 AddKeyXOR2_XORInst_4_0_U1 ( .A(MCOutput[16]), .B(SelectedKey[16]), 
        .Z(AddRoundKeyOutput[16]) );
  XOR2_X1 AddKeyXOR2_XORInst_4_1_U1 ( .A(MCOutput[17]), .B(SelectedKey[17]), 
        .Z(AddRoundKeyOutput[17]) );
  XOR2_X1 AddKeyXOR2_XORInst_4_2_U1 ( .A(MCOutput[18]), .B(SelectedKey[18]), 
        .Z(AddRoundKeyOutput[18]) );
  XOR2_X1 AddKeyXOR2_XORInst_4_3_U1 ( .A(MCOutput[19]), .B(SelectedKey[19]), 
        .Z(AddRoundKeyOutput[19]) );
  XOR2_X1 AddKeyXOR2_XORInst_5_0_U1 ( .A(MCOutput[20]), .B(SelectedKey[20]), 
        .Z(AddRoundKeyOutput[20]) );
  XOR2_X1 AddKeyXOR2_XORInst_5_1_U1 ( .A(MCOutput[21]), .B(SelectedKey[21]), 
        .Z(AddRoundKeyOutput[21]) );
  XOR2_X1 AddKeyXOR2_XORInst_5_2_U1 ( .A(MCOutput[22]), .B(SelectedKey[22]), 
        .Z(AddRoundKeyOutput[22]) );
  XOR2_X1 AddKeyXOR2_XORInst_5_3_U1 ( .A(MCOutput[23]), .B(SelectedKey[23]), 
        .Z(AddRoundKeyOutput[23]) );
  XOR2_X1 AddKeyXOR2_XORInst_6_0_U1 ( .A(MCOutput[24]), .B(SelectedKey[24]), 
        .Z(AddRoundKeyOutput[24]) );
  XOR2_X1 AddKeyXOR2_XORInst_6_1_U1 ( .A(MCOutput[25]), .B(SelectedKey[25]), 
        .Z(AddRoundKeyOutput[25]) );
  XOR2_X1 AddKeyXOR2_XORInst_6_2_U1 ( .A(MCOutput[26]), .B(SelectedKey[26]), 
        .Z(AddRoundKeyOutput[26]) );
  XOR2_X1 AddKeyXOR2_XORInst_6_3_U1 ( .A(MCOutput[27]), .B(SelectedKey[27]), 
        .Z(AddRoundKeyOutput[27]) );
  XOR2_X1 AddKeyXOR2_XORInst_7_0_U1 ( .A(MCOutput[28]), .B(SelectedKey[28]), 
        .Z(AddRoundKeyOutput[28]) );
  XOR2_X1 AddKeyXOR2_XORInst_7_1_U1 ( .A(MCOutput[29]), .B(SelectedKey[29]), 
        .Z(AddRoundKeyOutput[29]) );
  XOR2_X1 AddKeyXOR2_XORInst_7_2_U1 ( .A(MCOutput[30]), .B(SelectedKey[30]), 
        .Z(AddRoundKeyOutput[30]) );
  XOR2_X1 AddKeyXOR2_XORInst_7_3_U1 ( .A(MCOutput[31]), .B(SelectedKey[31]), 
        .Z(AddRoundKeyOutput[31]) );
  XOR2_X1 AddKeyXOR2_XORInst_8_0_U1 ( .A(MCOutput[32]), .B(SelectedKey[32]), 
        .Z(AddRoundKeyOutput[32]) );
  XOR2_X1 AddKeyXOR2_XORInst_8_1_U1 ( .A(MCOutput[33]), .B(SelectedKey[33]), 
        .Z(AddRoundKeyOutput[33]) );
  XOR2_X1 AddKeyXOR2_XORInst_8_2_U1 ( .A(MCOutput[34]), .B(SelectedKey[34]), 
        .Z(AddRoundKeyOutput[34]) );
  XOR2_X1 AddKeyXOR2_XORInst_8_3_U1 ( .A(MCOutput[35]), .B(SelectedKey[35]), 
        .Z(AddRoundKeyOutput[35]) );
  XOR2_X1 AddKeyXOR2_XORInst_9_0_U1 ( .A(MCOutput[36]), .B(SelectedKey[36]), 
        .Z(AddRoundKeyOutput[36]) );
  XOR2_X1 AddKeyXOR2_XORInst_9_1_U1 ( .A(MCOutput[37]), .B(SelectedKey[37]), 
        .Z(AddRoundKeyOutput[37]) );
  XOR2_X1 AddKeyXOR2_XORInst_9_2_U1 ( .A(MCOutput[38]), .B(SelectedKey[38]), 
        .Z(AddRoundKeyOutput[38]) );
  XOR2_X1 AddKeyXOR2_XORInst_9_3_U1 ( .A(MCOutput[39]), .B(SelectedKey[39]), 
        .Z(AddRoundKeyOutput[39]) );
  DFF_X1 StateReg_s_current_state_reg_0_ ( .D(AddRoundKeyOutput[0]), .CK(clk), 
        .Q(StateRegOutput[0]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_1_ ( .D(AddRoundKeyOutput[1]), .CK(clk), 
        .Q(StateRegOutput[1]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_2_ ( .D(AddRoundKeyOutput[2]), .CK(clk), 
        .Q(StateRegOutput[2]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_3_ ( .D(AddRoundKeyOutput[3]), .CK(clk), 
        .Q(StateRegOutput[3]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_4_ ( .D(AddRoundKeyOutput[4]), .CK(clk), 
        .Q(StateRegOutput[4]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_5_ ( .D(AddRoundKeyOutput[5]), .CK(clk), 
        .Q(StateRegOutput[5]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_6_ ( .D(AddRoundKeyOutput[6]), .CK(clk), 
        .Q(StateRegOutput[6]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_7_ ( .D(AddRoundKeyOutput[7]), .CK(clk), 
        .Q(StateRegOutput[7]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_8_ ( .D(AddRoundKeyOutput[8]), .CK(clk), 
        .Q(StateRegOutput[8]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_9_ ( .D(AddRoundKeyOutput[9]), .CK(clk), 
        .Q(StateRegOutput[9]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_10_ ( .D(AddRoundKeyOutput[10]), .CK(clk), .Q(StateRegOutput[10]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_11_ ( .D(AddRoundKeyOutput[11]), .CK(clk), .Q(StateRegOutput[11]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_12_ ( .D(AddRoundKeyOutput[12]), .CK(clk), .Q(StateRegOutput[12]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_13_ ( .D(AddRoundKeyOutput[13]), .CK(clk), .Q(StateRegOutput[13]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_14_ ( .D(AddRoundKeyOutput[14]), .CK(clk), .Q(StateRegOutput[14]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_15_ ( .D(AddRoundKeyOutput[15]), .CK(clk), .Q(StateRegOutput[15]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_16_ ( .D(AddRoundKeyOutput[16]), .CK(clk), .Q(StateRegOutput[16]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_17_ ( .D(AddRoundKeyOutput[17]), .CK(clk), .Q(StateRegOutput[17]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_18_ ( .D(AddRoundKeyOutput[18]), .CK(clk), .Q(StateRegOutput[18]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_19_ ( .D(AddRoundKeyOutput[19]), .CK(clk), .Q(StateRegOutput[19]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_20_ ( .D(AddRoundKeyOutput[20]), .CK(clk), .Q(StateRegOutput[20]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_21_ ( .D(AddRoundKeyOutput[21]), .CK(clk), .Q(StateRegOutput[21]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_22_ ( .D(AddRoundKeyOutput[22]), .CK(clk), .Q(StateRegOutput[22]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_23_ ( .D(AddRoundKeyOutput[23]), .CK(clk), .Q(StateRegOutput[23]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_24_ ( .D(AddRoundKeyOutput[24]), .CK(clk), .Q(StateRegOutput[24]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_25_ ( .D(AddRoundKeyOutput[25]), .CK(clk), .Q(StateRegOutput[25]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_26_ ( .D(AddRoundKeyOutput[26]), .CK(clk), .Q(StateRegOutput[26]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_27_ ( .D(AddRoundKeyOutput[27]), .CK(clk), .Q(StateRegOutput[27]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_28_ ( .D(AddRoundKeyOutput[28]), .CK(clk), .Q(StateRegOutput[28]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_29_ ( .D(AddRoundKeyOutput[29]), .CK(clk), .Q(StateRegOutput[29]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_30_ ( .D(AddRoundKeyOutput[30]), .CK(clk), .Q(StateRegOutput[30]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_31_ ( .D(AddRoundKeyOutput[31]), .CK(clk), .Q(StateRegOutput[31]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_32_ ( .D(AddRoundKeyOutput[32]), .CK(clk), .Q(StateRegOutput[32]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_33_ ( .D(AddRoundKeyOutput[33]), .CK(clk), .Q(StateRegOutput[33]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_34_ ( .D(AddRoundKeyOutput[34]), .CK(clk), .Q(StateRegOutput[34]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_35_ ( .D(AddRoundKeyOutput[35]), .CK(clk), .Q(StateRegOutput[35]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_36_ ( .D(AddRoundKeyOutput[36]), .CK(clk), .Q(StateRegOutput[36]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_37_ ( .D(AddRoundKeyOutput[37]), .CK(clk), .Q(StateRegOutput[37]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_38_ ( .D(AddRoundKeyOutput[38]), .CK(clk), .Q(StateRegOutput[38]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_39_ ( .D(AddRoundKeyOutput[39]), .CK(clk), .Q(StateRegOutput[39]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_40_ ( .D(AddRoundKeyOutput[40]), .CK(clk), .Q(StateRegOutput[40]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_41_ ( .D(AddRoundKeyOutput[41]), .CK(clk), .Q(StateRegOutput[41]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_42_ ( .D(AddRoundKeyOutput[42]), .CK(clk), .Q(StateRegOutput[42]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_43_ ( .D(AddRoundKeyOutput[43]), .CK(clk), .Q(StateRegOutput[43]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_44_ ( .D(AddRoundKeyOutput[44]), .CK(clk), .Q(StateRegOutput[44]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_45_ ( .D(AddRoundKeyOutput[45]), .CK(clk), .Q(StateRegOutput[45]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_46_ ( .D(AddRoundKeyOutput[46]), .CK(clk), .Q(StateRegOutput[46]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_47_ ( .D(AddRoundKeyOutput[47]), .CK(clk), .Q(StateRegOutput[47]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_48_ ( .D(AddRoundKeyOutput[48]), .CK(clk), .Q(StateRegOutput[48]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_49_ ( .D(AddRoundKeyOutput[49]), .CK(clk), .Q(StateRegOutput[49]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_50_ ( .D(AddRoundKeyOutput[50]), .CK(clk), .Q(StateRegOutput[50]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_51_ ( .D(AddRoundKeyOutput[51]), .CK(clk), .Q(StateRegOutput[51]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_52_ ( .D(AddRoundKeyOutput[52]), .CK(clk), .Q(StateRegOutput[52]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_53_ ( .D(AddRoundKeyOutput[53]), .CK(clk), .Q(StateRegOutput[53]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_54_ ( .D(AddRoundKeyOutput[54]), .CK(clk), .Q(StateRegOutput[54]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_55_ ( .D(AddRoundKeyOutput[55]), .CK(clk), .Q(StateRegOutput[55]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_56_ ( .D(AddRoundKeyOutput[56]), .CK(clk), .Q(StateRegOutput[56]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_57_ ( .D(AddRoundKeyOutput[57]), .CK(clk), .Q(StateRegOutput[57]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_58_ ( .D(AddRoundKeyOutput[58]), .CK(clk), .Q(StateRegOutput[58]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_59_ ( .D(AddRoundKeyOutput[59]), .CK(clk), .Q(StateRegOutput[59]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_60_ ( .D(AddRoundKeyOutput[60]), .CK(clk), .Q(StateRegOutput[60]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_61_ ( .D(AddRoundKeyOutput[61]), .CK(clk), .Q(StateRegOutput[61]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_62_ ( .D(AddRoundKeyOutput[62]), .CK(clk), .Q(StateRegOutput[62]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_63_ ( .D(AddRoundKeyOutput[63]), .CK(clk), .Q(StateRegOutput[63]), .QN() );
  XNOR2_X1 F_StateRegOutput_Inst_LFInst_0_LFInst_0_U2 ( .A(
        F_StateRegOutput_Inst_LFInst_0_LFInst_0_n3), .B(StateRegOutput[2]), 
        .ZN(StateRegOutputF[0]) );
  XNOR2_X1 F_StateRegOutput_Inst_LFInst_0_LFInst_0_U1 ( .A(StateRegOutput[0]), 
        .B(StateRegOutput[1]), .ZN(F_StateRegOutput_Inst_LFInst_0_LFInst_0_n3)
         );
  XNOR2_X1 F_StateRegOutput_Inst_LFInst_0_LFInst_1_U2 ( .A(
        F_StateRegOutput_Inst_LFInst_0_LFInst_1_n3), .B(StateRegOutput[3]), 
        .ZN(StateRegOutputF[1]) );
  XNOR2_X1 F_StateRegOutput_Inst_LFInst_0_LFInst_1_U1 ( .A(StateRegOutput[0]), 
        .B(StateRegOutput[1]), .ZN(F_StateRegOutput_Inst_LFInst_0_LFInst_1_n3)
         );
  XOR2_X1 F_StateRegOutput_Inst_LFInst_0_LFInst_2_U1 ( .A(StateRegOutput[0]), 
        .B(StateRegOutput[2]), .Z(StateRegOutputF[2]) );
  XOR2_X1 F_StateRegOutput_Inst_LFInst_0_LFInst_3_U1 ( .A(StateRegOutput[0]), 
        .B(StateRegOutput[3]), .Z(StateRegOutputF[3]) );
  XOR2_X1 F_StateRegOutput_Inst_LFInst_0_LFInst_4_U1 ( .A(StateRegOutput[1]), 
        .B(StateRegOutput[2]), .Z(StateRegOutputF[4]) );
  XOR2_X1 F_StateRegOutput_Inst_LFInst_0_LFInst_5_U1 ( .A(StateRegOutput[1]), 
        .B(StateRegOutput[3]), .Z(StateRegOutputF[5]) );
  XOR2_X1 F_StateRegOutput_Inst_LFInst_0_LFInst_6_U1 ( .A(StateRegOutput[2]), 
        .B(StateRegOutput[3]), .Z(StateRegOutputF[6]) );
  XNOR2_X1 F_StateRegOutput_Inst_LFInst_1_LFInst_0_U2 ( .A(
        F_StateRegOutput_Inst_LFInst_1_LFInst_0_n3), .B(StateRegOutput[6]), 
        .ZN(StateRegOutputF[7]) );
  XNOR2_X1 F_StateRegOutput_Inst_LFInst_1_LFInst_0_U1 ( .A(StateRegOutput[4]), 
        .B(StateRegOutput[5]), .ZN(F_StateRegOutput_Inst_LFInst_1_LFInst_0_n3)
         );
  XNOR2_X1 F_StateRegOutput_Inst_LFInst_1_LFInst_1_U2 ( .A(
        F_StateRegOutput_Inst_LFInst_1_LFInst_1_n3), .B(StateRegOutput[7]), 
        .ZN(StateRegOutputF[8]) );
  XNOR2_X1 F_StateRegOutput_Inst_LFInst_1_LFInst_1_U1 ( .A(StateRegOutput[4]), 
        .B(StateRegOutput[5]), .ZN(F_StateRegOutput_Inst_LFInst_1_LFInst_1_n3)
         );
  XOR2_X1 F_StateRegOutput_Inst_LFInst_1_LFInst_2_U1 ( .A(StateRegOutput[4]), 
        .B(StateRegOutput[6]), .Z(StateRegOutputF[9]) );
  XOR2_X1 F_StateRegOutput_Inst_LFInst_1_LFInst_3_U1 ( .A(StateRegOutput[4]), 
        .B(StateRegOutput[7]), .Z(StateRegOutputF[10]) );
  XOR2_X1 F_StateRegOutput_Inst_LFInst_1_LFInst_4_U1 ( .A(StateRegOutput[5]), 
        .B(StateRegOutput[6]), .Z(StateRegOutputF[11]) );
  XOR2_X1 F_StateRegOutput_Inst_LFInst_1_LFInst_5_U1 ( .A(StateRegOutput[5]), 
        .B(StateRegOutput[7]), .Z(StateRegOutputF[12]) );
  XOR2_X1 F_StateRegOutput_Inst_LFInst_1_LFInst_6_U1 ( .A(StateRegOutput[6]), 
        .B(StateRegOutput[7]), .Z(StateRegOutputF[13]) );
  XNOR2_X1 F_StateRegOutput_Inst_LFInst_2_LFInst_0_U2 ( .A(
        F_StateRegOutput_Inst_LFInst_2_LFInst_0_n3), .B(StateRegOutput[10]), 
        .ZN(StateRegOutputF[14]) );
  XNOR2_X1 F_StateRegOutput_Inst_LFInst_2_LFInst_0_U1 ( .A(StateRegOutput[8]), 
        .B(StateRegOutput[9]), .ZN(F_StateRegOutput_Inst_LFInst_2_LFInst_0_n3)
         );
  XNOR2_X1 F_StateRegOutput_Inst_LFInst_2_LFInst_1_U2 ( .A(
        F_StateRegOutput_Inst_LFInst_2_LFInst_1_n3), .B(StateRegOutput[11]), 
        .ZN(StateRegOutputF[15]) );
  XNOR2_X1 F_StateRegOutput_Inst_LFInst_2_LFInst_1_U1 ( .A(StateRegOutput[8]), 
        .B(StateRegOutput[9]), .ZN(F_StateRegOutput_Inst_LFInst_2_LFInst_1_n3)
         );
  XOR2_X1 F_StateRegOutput_Inst_LFInst_2_LFInst_2_U1 ( .A(StateRegOutput[8]), 
        .B(StateRegOutput[10]), .Z(StateRegOutputF[16]) );
  XOR2_X1 F_StateRegOutput_Inst_LFInst_2_LFInst_3_U1 ( .A(StateRegOutput[8]), 
        .B(StateRegOutput[11]), .Z(StateRegOutputF[17]) );
  XOR2_X1 F_StateRegOutput_Inst_LFInst_2_LFInst_4_U1 ( .A(StateRegOutput[9]), 
        .B(StateRegOutput[10]), .Z(StateRegOutputF[18]) );
  XOR2_X1 F_StateRegOutput_Inst_LFInst_2_LFInst_5_U1 ( .A(StateRegOutput[9]), 
        .B(StateRegOutput[11]), .Z(StateRegOutputF[19]) );
  XOR2_X1 F_StateRegOutput_Inst_LFInst_2_LFInst_6_U1 ( .A(StateRegOutput[10]), 
        .B(StateRegOutput[11]), .Z(StateRegOutputF[20]) );
  XNOR2_X1 F_StateRegOutput_Inst_LFInst_3_LFInst_0_U2 ( .A(
        F_StateRegOutput_Inst_LFInst_3_LFInst_0_n3), .B(StateRegOutput[14]), 
        .ZN(StateRegOutputF[21]) );
  XNOR2_X1 F_StateRegOutput_Inst_LFInst_3_LFInst_0_U1 ( .A(StateRegOutput[12]), 
        .B(StateRegOutput[13]), .ZN(F_StateRegOutput_Inst_LFInst_3_LFInst_0_n3) );
  XNOR2_X1 F_StateRegOutput_Inst_LFInst_3_LFInst_1_U2 ( .A(
        F_StateRegOutput_Inst_LFInst_3_LFInst_1_n3), .B(StateRegOutput[15]), 
        .ZN(StateRegOutputF[22]) );
  XNOR2_X1 F_StateRegOutput_Inst_LFInst_3_LFInst_1_U1 ( .A(StateRegOutput[12]), 
        .B(StateRegOutput[13]), .ZN(F_StateRegOutput_Inst_LFInst_3_LFInst_1_n3) );
  XOR2_X1 F_StateRegOutput_Inst_LFInst_3_LFInst_2_U1 ( .A(StateRegOutput[12]), 
        .B(StateRegOutput[14]), .Z(StateRegOutputF[23]) );
  XOR2_X1 F_StateRegOutput_Inst_LFInst_3_LFInst_3_U1 ( .A(StateRegOutput[12]), 
        .B(StateRegOutput[15]), .Z(StateRegOutputF[24]) );
  XOR2_X1 F_StateRegOutput_Inst_LFInst_3_LFInst_4_U1 ( .A(StateRegOutput[13]), 
        .B(StateRegOutput[14]), .Z(StateRegOutputF[25]) );
  XOR2_X1 F_StateRegOutput_Inst_LFInst_3_LFInst_5_U1 ( .A(StateRegOutput[13]), 
        .B(StateRegOutput[15]), .Z(StateRegOutputF[26]) );
  XOR2_X1 F_StateRegOutput_Inst_LFInst_3_LFInst_6_U1 ( .A(StateRegOutput[14]), 
        .B(StateRegOutput[15]), .Z(StateRegOutputF[27]) );
  XNOR2_X1 F_StateRegOutput_Inst_LFInst_4_LFInst_0_U2 ( .A(
        F_StateRegOutput_Inst_LFInst_4_LFInst_0_n3), .B(StateRegOutput[18]), 
        .ZN(StateRegOutputF[28]) );
  XNOR2_X1 F_StateRegOutput_Inst_LFInst_4_LFInst_0_U1 ( .A(StateRegOutput[16]), 
        .B(StateRegOutput[17]), .ZN(F_StateRegOutput_Inst_LFInst_4_LFInst_0_n3) );
  XNOR2_X1 F_StateRegOutput_Inst_LFInst_4_LFInst_1_U2 ( .A(
        F_StateRegOutput_Inst_LFInst_4_LFInst_1_n3), .B(StateRegOutput[19]), 
        .ZN(StateRegOutputF[29]) );
  XNOR2_X1 F_StateRegOutput_Inst_LFInst_4_LFInst_1_U1 ( .A(StateRegOutput[16]), 
        .B(StateRegOutput[17]), .ZN(F_StateRegOutput_Inst_LFInst_4_LFInst_1_n3) );
  XOR2_X1 F_StateRegOutput_Inst_LFInst_4_LFInst_2_U1 ( .A(StateRegOutput[16]), 
        .B(StateRegOutput[18]), .Z(StateRegOutputF[30]) );
  XOR2_X1 F_StateRegOutput_Inst_LFInst_4_LFInst_3_U1 ( .A(StateRegOutput[16]), 
        .B(StateRegOutput[19]), .Z(StateRegOutputF[31]) );
  XOR2_X1 F_StateRegOutput_Inst_LFInst_4_LFInst_4_U1 ( .A(StateRegOutput[17]), 
        .B(StateRegOutput[18]), .Z(StateRegOutputF[32]) );
  XOR2_X1 F_StateRegOutput_Inst_LFInst_4_LFInst_5_U1 ( .A(StateRegOutput[17]), 
        .B(StateRegOutput[19]), .Z(StateRegOutputF[33]) );
  XOR2_X1 F_StateRegOutput_Inst_LFInst_4_LFInst_6_U1 ( .A(StateRegOutput[18]), 
        .B(StateRegOutput[19]), .Z(StateRegOutputF[34]) );
  XNOR2_X1 F_StateRegOutput_Inst_LFInst_5_LFInst_0_U2 ( .A(
        F_StateRegOutput_Inst_LFInst_5_LFInst_0_n3), .B(StateRegOutput[22]), 
        .ZN(StateRegOutputF[35]) );
  XNOR2_X1 F_StateRegOutput_Inst_LFInst_5_LFInst_0_U1 ( .A(StateRegOutput[20]), 
        .B(StateRegOutput[21]), .ZN(F_StateRegOutput_Inst_LFInst_5_LFInst_0_n3) );
  XNOR2_X1 F_StateRegOutput_Inst_LFInst_5_LFInst_1_U2 ( .A(
        F_StateRegOutput_Inst_LFInst_5_LFInst_1_n3), .B(StateRegOutput[23]), 
        .ZN(StateRegOutputF[36]) );
  XNOR2_X1 F_StateRegOutput_Inst_LFInst_5_LFInst_1_U1 ( .A(StateRegOutput[20]), 
        .B(StateRegOutput[21]), .ZN(F_StateRegOutput_Inst_LFInst_5_LFInst_1_n3) );
  XOR2_X1 F_StateRegOutput_Inst_LFInst_5_LFInst_2_U1 ( .A(StateRegOutput[20]), 
        .B(StateRegOutput[22]), .Z(StateRegOutputF[37]) );
  XOR2_X1 F_StateRegOutput_Inst_LFInst_5_LFInst_3_U1 ( .A(StateRegOutput[20]), 
        .B(StateRegOutput[23]), .Z(StateRegOutputF[38]) );
  XOR2_X1 F_StateRegOutput_Inst_LFInst_5_LFInst_4_U1 ( .A(StateRegOutput[21]), 
        .B(StateRegOutput[22]), .Z(StateRegOutputF[39]) );
  XOR2_X1 F_StateRegOutput_Inst_LFInst_5_LFInst_5_U1 ( .A(StateRegOutput[21]), 
        .B(StateRegOutput[23]), .Z(StateRegOutputF[40]) );
  XOR2_X1 F_StateRegOutput_Inst_LFInst_5_LFInst_6_U1 ( .A(StateRegOutput[22]), 
        .B(StateRegOutput[23]), .Z(StateRegOutputF[41]) );
  XNOR2_X1 F_StateRegOutput_Inst_LFInst_6_LFInst_0_U2 ( .A(
        F_StateRegOutput_Inst_LFInst_6_LFInst_0_n3), .B(StateRegOutput[26]), 
        .ZN(StateRegOutputF[42]) );
  XNOR2_X1 F_StateRegOutput_Inst_LFInst_6_LFInst_0_U1 ( .A(StateRegOutput[24]), 
        .B(StateRegOutput[25]), .ZN(F_StateRegOutput_Inst_LFInst_6_LFInst_0_n3) );
  XNOR2_X1 F_StateRegOutput_Inst_LFInst_6_LFInst_1_U2 ( .A(
        F_StateRegOutput_Inst_LFInst_6_LFInst_1_n3), .B(StateRegOutput[27]), 
        .ZN(StateRegOutputF[43]) );
  XNOR2_X1 F_StateRegOutput_Inst_LFInst_6_LFInst_1_U1 ( .A(StateRegOutput[24]), 
        .B(StateRegOutput[25]), .ZN(F_StateRegOutput_Inst_LFInst_6_LFInst_1_n3) );
  XOR2_X1 F_StateRegOutput_Inst_LFInst_6_LFInst_2_U1 ( .A(StateRegOutput[24]), 
        .B(StateRegOutput[26]), .Z(StateRegOutputF[44]) );
  XOR2_X1 F_StateRegOutput_Inst_LFInst_6_LFInst_3_U1 ( .A(StateRegOutput[24]), 
        .B(StateRegOutput[27]), .Z(StateRegOutputF[45]) );
  XOR2_X1 F_StateRegOutput_Inst_LFInst_6_LFInst_4_U1 ( .A(StateRegOutput[25]), 
        .B(StateRegOutput[26]), .Z(StateRegOutputF[46]) );
  XOR2_X1 F_StateRegOutput_Inst_LFInst_6_LFInst_5_U1 ( .A(StateRegOutput[25]), 
        .B(StateRegOutput[27]), .Z(StateRegOutputF[47]) );
  XOR2_X1 F_StateRegOutput_Inst_LFInst_6_LFInst_6_U1 ( .A(StateRegOutput[26]), 
        .B(StateRegOutput[27]), .Z(StateRegOutputF[48]) );
  XNOR2_X1 F_StateRegOutput_Inst_LFInst_7_LFInst_0_U2 ( .A(
        F_StateRegOutput_Inst_LFInst_7_LFInst_0_n3), .B(StateRegOutput[30]), 
        .ZN(StateRegOutputF[49]) );
  XNOR2_X1 F_StateRegOutput_Inst_LFInst_7_LFInst_0_U1 ( .A(StateRegOutput[28]), 
        .B(StateRegOutput[29]), .ZN(F_StateRegOutput_Inst_LFInst_7_LFInst_0_n3) );
  XNOR2_X1 F_StateRegOutput_Inst_LFInst_7_LFInst_1_U2 ( .A(
        F_StateRegOutput_Inst_LFInst_7_LFInst_1_n3), .B(StateRegOutput[31]), 
        .ZN(StateRegOutputF[50]) );
  XNOR2_X1 F_StateRegOutput_Inst_LFInst_7_LFInst_1_U1 ( .A(StateRegOutput[28]), 
        .B(StateRegOutput[29]), .ZN(F_StateRegOutput_Inst_LFInst_7_LFInst_1_n3) );
  XOR2_X1 F_StateRegOutput_Inst_LFInst_7_LFInst_2_U1 ( .A(StateRegOutput[28]), 
        .B(StateRegOutput[30]), .Z(StateRegOutputF[51]) );
  XOR2_X1 F_StateRegOutput_Inst_LFInst_7_LFInst_3_U1 ( .A(StateRegOutput[28]), 
        .B(StateRegOutput[31]), .Z(StateRegOutputF[52]) );
  XOR2_X1 F_StateRegOutput_Inst_LFInst_7_LFInst_4_U1 ( .A(StateRegOutput[29]), 
        .B(StateRegOutput[30]), .Z(StateRegOutputF[53]) );
  XOR2_X1 F_StateRegOutput_Inst_LFInst_7_LFInst_5_U1 ( .A(StateRegOutput[29]), 
        .B(StateRegOutput[31]), .Z(StateRegOutputF[54]) );
  XOR2_X1 F_StateRegOutput_Inst_LFInst_7_LFInst_6_U1 ( .A(StateRegOutput[30]), 
        .B(StateRegOutput[31]), .Z(StateRegOutputF[55]) );
  XNOR2_X1 F_StateRegOutput_Inst_LFInst_8_LFInst_0_U2 ( .A(
        F_StateRegOutput_Inst_LFInst_8_LFInst_0_n3), .B(StateRegOutput[34]), 
        .ZN(StateRegOutputF[56]) );
  XNOR2_X1 F_StateRegOutput_Inst_LFInst_8_LFInst_0_U1 ( .A(StateRegOutput[32]), 
        .B(StateRegOutput[33]), .ZN(F_StateRegOutput_Inst_LFInst_8_LFInst_0_n3) );
  XNOR2_X1 F_StateRegOutput_Inst_LFInst_8_LFInst_1_U2 ( .A(
        F_StateRegOutput_Inst_LFInst_8_LFInst_1_n3), .B(StateRegOutput[35]), 
        .ZN(StateRegOutputF[57]) );
  XNOR2_X1 F_StateRegOutput_Inst_LFInst_8_LFInst_1_U1 ( .A(StateRegOutput[32]), 
        .B(StateRegOutput[33]), .ZN(F_StateRegOutput_Inst_LFInst_8_LFInst_1_n3) );
  XOR2_X1 F_StateRegOutput_Inst_LFInst_8_LFInst_2_U1 ( .A(StateRegOutput[32]), 
        .B(StateRegOutput[34]), .Z(StateRegOutputF[58]) );
  XOR2_X1 F_StateRegOutput_Inst_LFInst_8_LFInst_3_U1 ( .A(StateRegOutput[32]), 
        .B(StateRegOutput[35]), .Z(StateRegOutputF[59]) );
  XOR2_X1 F_StateRegOutput_Inst_LFInst_8_LFInst_4_U1 ( .A(StateRegOutput[33]), 
        .B(StateRegOutput[34]), .Z(StateRegOutputF[60]) );
  XOR2_X1 F_StateRegOutput_Inst_LFInst_8_LFInst_5_U1 ( .A(StateRegOutput[33]), 
        .B(StateRegOutput[35]), .Z(StateRegOutputF[61]) );
  XOR2_X1 F_StateRegOutput_Inst_LFInst_8_LFInst_6_U1 ( .A(StateRegOutput[34]), 
        .B(StateRegOutput[35]), .Z(StateRegOutputF[62]) );
  XNOR2_X1 F_StateRegOutput_Inst_LFInst_9_LFInst_0_U2 ( .A(
        F_StateRegOutput_Inst_LFInst_9_LFInst_0_n3), .B(StateRegOutput[38]), 
        .ZN(StateRegOutputF[63]) );
  XNOR2_X1 F_StateRegOutput_Inst_LFInst_9_LFInst_0_U1 ( .A(StateRegOutput[36]), 
        .B(StateRegOutput[37]), .ZN(F_StateRegOutput_Inst_LFInst_9_LFInst_0_n3) );
  XNOR2_X1 F_StateRegOutput_Inst_LFInst_9_LFInst_1_U2 ( .A(
        F_StateRegOutput_Inst_LFInst_9_LFInst_1_n3), .B(StateRegOutput[39]), 
        .ZN(StateRegOutputF[64]) );
  XNOR2_X1 F_StateRegOutput_Inst_LFInst_9_LFInst_1_U1 ( .A(StateRegOutput[36]), 
        .B(StateRegOutput[37]), .ZN(F_StateRegOutput_Inst_LFInst_9_LFInst_1_n3) );
  XOR2_X1 F_StateRegOutput_Inst_LFInst_9_LFInst_2_U1 ( .A(StateRegOutput[36]), 
        .B(StateRegOutput[38]), .Z(StateRegOutputF[65]) );
  XOR2_X1 F_StateRegOutput_Inst_LFInst_9_LFInst_3_U1 ( .A(StateRegOutput[36]), 
        .B(StateRegOutput[39]), .Z(StateRegOutputF[66]) );
  XOR2_X1 F_StateRegOutput_Inst_LFInst_9_LFInst_4_U1 ( .A(StateRegOutput[37]), 
        .B(StateRegOutput[38]), .Z(StateRegOutputF[67]) );
  XOR2_X1 F_StateRegOutput_Inst_LFInst_9_LFInst_5_U1 ( .A(StateRegOutput[37]), 
        .B(StateRegOutput[39]), .Z(StateRegOutputF[68]) );
  XOR2_X1 F_StateRegOutput_Inst_LFInst_9_LFInst_6_U1 ( .A(StateRegOutput[38]), 
        .B(StateRegOutput[39]), .Z(StateRegOutputF[69]) );
  XNOR2_X1 F_StateRegOutput_Inst_LFInst_10_LFInst_0_U2 ( .A(
        F_StateRegOutput_Inst_LFInst_10_LFInst_0_n3), .B(StateRegOutput[42]), 
        .ZN(StateRegOutputF[70]) );
  XNOR2_X1 F_StateRegOutput_Inst_LFInst_10_LFInst_0_U1 ( .A(StateRegOutput[40]), .B(StateRegOutput[41]), .ZN(F_StateRegOutput_Inst_LFInst_10_LFInst_0_n3) );
  XNOR2_X1 F_StateRegOutput_Inst_LFInst_10_LFInst_1_U2 ( .A(
        F_StateRegOutput_Inst_LFInst_10_LFInst_1_n3), .B(StateRegOutput[43]), 
        .ZN(StateRegOutputF[71]) );
  XNOR2_X1 F_StateRegOutput_Inst_LFInst_10_LFInst_1_U1 ( .A(StateRegOutput[40]), .B(StateRegOutput[41]), .ZN(F_StateRegOutput_Inst_LFInst_10_LFInst_1_n3) );
  XOR2_X1 F_StateRegOutput_Inst_LFInst_10_LFInst_2_U1 ( .A(StateRegOutput[40]), 
        .B(StateRegOutput[42]), .Z(StateRegOutputF[72]) );
  XOR2_X1 F_StateRegOutput_Inst_LFInst_10_LFInst_3_U1 ( .A(StateRegOutput[40]), 
        .B(StateRegOutput[43]), .Z(StateRegOutputF[73]) );
  XOR2_X1 F_StateRegOutput_Inst_LFInst_10_LFInst_4_U1 ( .A(StateRegOutput[41]), 
        .B(StateRegOutput[42]), .Z(StateRegOutputF[74]) );
  XOR2_X1 F_StateRegOutput_Inst_LFInst_10_LFInst_5_U1 ( .A(StateRegOutput[41]), 
        .B(StateRegOutput[43]), .Z(StateRegOutputF[75]) );
  XOR2_X1 F_StateRegOutput_Inst_LFInst_10_LFInst_6_U1 ( .A(StateRegOutput[42]), 
        .B(StateRegOutput[43]), .Z(StateRegOutputF[76]) );
  XNOR2_X1 F_StateRegOutput_Inst_LFInst_11_LFInst_0_U2 ( .A(
        F_StateRegOutput_Inst_LFInst_11_LFInst_0_n3), .B(StateRegOutput[46]), 
        .ZN(StateRegOutputF[77]) );
  XNOR2_X1 F_StateRegOutput_Inst_LFInst_11_LFInst_0_U1 ( .A(StateRegOutput[44]), .B(StateRegOutput[45]), .ZN(F_StateRegOutput_Inst_LFInst_11_LFInst_0_n3) );
  XNOR2_X1 F_StateRegOutput_Inst_LFInst_11_LFInst_1_U2 ( .A(
        F_StateRegOutput_Inst_LFInst_11_LFInst_1_n3), .B(StateRegOutput[47]), 
        .ZN(StateRegOutputF[78]) );
  XNOR2_X1 F_StateRegOutput_Inst_LFInst_11_LFInst_1_U1 ( .A(StateRegOutput[44]), .B(StateRegOutput[45]), .ZN(F_StateRegOutput_Inst_LFInst_11_LFInst_1_n3) );
  XOR2_X1 F_StateRegOutput_Inst_LFInst_11_LFInst_2_U1 ( .A(StateRegOutput[44]), 
        .B(StateRegOutput[46]), .Z(StateRegOutputF[79]) );
  XOR2_X1 F_StateRegOutput_Inst_LFInst_11_LFInst_3_U1 ( .A(StateRegOutput[44]), 
        .B(StateRegOutput[47]), .Z(StateRegOutputF[80]) );
  XOR2_X1 F_StateRegOutput_Inst_LFInst_11_LFInst_4_U1 ( .A(StateRegOutput[45]), 
        .B(StateRegOutput[46]), .Z(StateRegOutputF[81]) );
  XOR2_X1 F_StateRegOutput_Inst_LFInst_11_LFInst_5_U1 ( .A(StateRegOutput[45]), 
        .B(StateRegOutput[47]), .Z(StateRegOutputF[82]) );
  XOR2_X1 F_StateRegOutput_Inst_LFInst_11_LFInst_6_U1 ( .A(StateRegOutput[46]), 
        .B(StateRegOutput[47]), .Z(StateRegOutputF[83]) );
  XNOR2_X1 F_StateRegOutput_Inst_LFInst_12_LFInst_0_U2 ( .A(
        F_StateRegOutput_Inst_LFInst_12_LFInst_0_n3), .B(StateRegOutput[50]), 
        .ZN(StateRegOutputF[84]) );
  XNOR2_X1 F_StateRegOutput_Inst_LFInst_12_LFInst_0_U1 ( .A(StateRegOutput[48]), .B(StateRegOutput[49]), .ZN(F_StateRegOutput_Inst_LFInst_12_LFInst_0_n3) );
  XNOR2_X1 F_StateRegOutput_Inst_LFInst_12_LFInst_1_U2 ( .A(
        F_StateRegOutput_Inst_LFInst_12_LFInst_1_n3), .B(StateRegOutput[51]), 
        .ZN(StateRegOutputF[85]) );
  XNOR2_X1 F_StateRegOutput_Inst_LFInst_12_LFInst_1_U1 ( .A(StateRegOutput[48]), .B(StateRegOutput[49]), .ZN(F_StateRegOutput_Inst_LFInst_12_LFInst_1_n3) );
  XOR2_X1 F_StateRegOutput_Inst_LFInst_12_LFInst_2_U1 ( .A(StateRegOutput[48]), 
        .B(StateRegOutput[50]), .Z(StateRegOutputF[86]) );
  XOR2_X1 F_StateRegOutput_Inst_LFInst_12_LFInst_3_U1 ( .A(StateRegOutput[48]), 
        .B(StateRegOutput[51]), .Z(StateRegOutputF[87]) );
  XOR2_X1 F_StateRegOutput_Inst_LFInst_12_LFInst_4_U1 ( .A(StateRegOutput[49]), 
        .B(StateRegOutput[50]), .Z(StateRegOutputF[88]) );
  XOR2_X1 F_StateRegOutput_Inst_LFInst_12_LFInst_5_U1 ( .A(StateRegOutput[49]), 
        .B(StateRegOutput[51]), .Z(StateRegOutputF[89]) );
  XOR2_X1 F_StateRegOutput_Inst_LFInst_12_LFInst_6_U1 ( .A(StateRegOutput[50]), 
        .B(StateRegOutput[51]), .Z(StateRegOutputF[90]) );
  XNOR2_X1 F_StateRegOutput_Inst_LFInst_13_LFInst_0_U2 ( .A(
        F_StateRegOutput_Inst_LFInst_13_LFInst_0_n3), .B(StateRegOutput[54]), 
        .ZN(StateRegOutputF[91]) );
  XNOR2_X1 F_StateRegOutput_Inst_LFInst_13_LFInst_0_U1 ( .A(StateRegOutput[52]), .B(StateRegOutput[53]), .ZN(F_StateRegOutput_Inst_LFInst_13_LFInst_0_n3) );
  XNOR2_X1 F_StateRegOutput_Inst_LFInst_13_LFInst_1_U2 ( .A(
        F_StateRegOutput_Inst_LFInst_13_LFInst_1_n3), .B(StateRegOutput[55]), 
        .ZN(StateRegOutputF[92]) );
  XNOR2_X1 F_StateRegOutput_Inst_LFInst_13_LFInst_1_U1 ( .A(StateRegOutput[52]), .B(StateRegOutput[53]), .ZN(F_StateRegOutput_Inst_LFInst_13_LFInst_1_n3) );
  XOR2_X1 F_StateRegOutput_Inst_LFInst_13_LFInst_2_U1 ( .A(StateRegOutput[52]), 
        .B(StateRegOutput[54]), .Z(StateRegOutputF[93]) );
  XOR2_X1 F_StateRegOutput_Inst_LFInst_13_LFInst_3_U1 ( .A(StateRegOutput[52]), 
        .B(StateRegOutput[55]), .Z(StateRegOutputF[94]) );
  XOR2_X1 F_StateRegOutput_Inst_LFInst_13_LFInst_4_U1 ( .A(StateRegOutput[53]), 
        .B(StateRegOutput[54]), .Z(StateRegOutputF[95]) );
  XOR2_X1 F_StateRegOutput_Inst_LFInst_13_LFInst_5_U1 ( .A(StateRegOutput[53]), 
        .B(StateRegOutput[55]), .Z(StateRegOutputF[96]) );
  XOR2_X1 F_StateRegOutput_Inst_LFInst_13_LFInst_6_U1 ( .A(StateRegOutput[54]), 
        .B(StateRegOutput[55]), .Z(StateRegOutputF[97]) );
  XNOR2_X1 F_StateRegOutput_Inst_LFInst_14_LFInst_0_U2 ( .A(
        F_StateRegOutput_Inst_LFInst_14_LFInst_0_n3), .B(StateRegOutput[58]), 
        .ZN(StateRegOutputF[98]) );
  XNOR2_X1 F_StateRegOutput_Inst_LFInst_14_LFInst_0_U1 ( .A(StateRegOutput[56]), .B(StateRegOutput[57]), .ZN(F_StateRegOutput_Inst_LFInst_14_LFInst_0_n3) );
  XNOR2_X1 F_StateRegOutput_Inst_LFInst_14_LFInst_1_U2 ( .A(
        F_StateRegOutput_Inst_LFInst_14_LFInst_1_n3), .B(StateRegOutput[59]), 
        .ZN(StateRegOutputF[99]) );
  XNOR2_X1 F_StateRegOutput_Inst_LFInst_14_LFInst_1_U1 ( .A(StateRegOutput[56]), .B(StateRegOutput[57]), .ZN(F_StateRegOutput_Inst_LFInst_14_LFInst_1_n3) );
  XOR2_X1 F_StateRegOutput_Inst_LFInst_14_LFInst_2_U1 ( .A(StateRegOutput[56]), 
        .B(StateRegOutput[58]), .Z(StateRegOutputF[100]) );
  XOR2_X1 F_StateRegOutput_Inst_LFInst_14_LFInst_3_U1 ( .A(StateRegOutput[56]), 
        .B(StateRegOutput[59]), .Z(StateRegOutputF[101]) );
  XOR2_X1 F_StateRegOutput_Inst_LFInst_14_LFInst_4_U1 ( .A(StateRegOutput[57]), 
        .B(StateRegOutput[58]), .Z(StateRegOutputF[102]) );
  XOR2_X1 F_StateRegOutput_Inst_LFInst_14_LFInst_5_U1 ( .A(StateRegOutput[57]), 
        .B(StateRegOutput[59]), .Z(StateRegOutputF[103]) );
  XOR2_X1 F_StateRegOutput_Inst_LFInst_14_LFInst_6_U1 ( .A(StateRegOutput[58]), 
        .B(StateRegOutput[59]), .Z(StateRegOutputF[104]) );
  XNOR2_X1 F_StateRegOutput_Inst_LFInst_15_LFInst_0_U2 ( .A(
        F_StateRegOutput_Inst_LFInst_15_LFInst_0_n3), .B(StateRegOutput[62]), 
        .ZN(StateRegOutputF[105]) );
  XNOR2_X1 F_StateRegOutput_Inst_LFInst_15_LFInst_0_U1 ( .A(StateRegOutput[60]), .B(StateRegOutput[61]), .ZN(F_StateRegOutput_Inst_LFInst_15_LFInst_0_n3) );
  XNOR2_X1 F_StateRegOutput_Inst_LFInst_15_LFInst_1_U2 ( .A(
        F_StateRegOutput_Inst_LFInst_15_LFInst_1_n3), .B(StateRegOutput[63]), 
        .ZN(StateRegOutputF[106]) );
  XNOR2_X1 F_StateRegOutput_Inst_LFInst_15_LFInst_1_U1 ( .A(StateRegOutput[60]), .B(StateRegOutput[61]), .ZN(F_StateRegOutput_Inst_LFInst_15_LFInst_1_n3) );
  XOR2_X1 F_StateRegOutput_Inst_LFInst_15_LFInst_2_U1 ( .A(StateRegOutput[60]), 
        .B(StateRegOutput[62]), .Z(StateRegOutputF[107]) );
  XOR2_X1 F_StateRegOutput_Inst_LFInst_15_LFInst_3_U1 ( .A(StateRegOutput[60]), 
        .B(StateRegOutput[63]), .Z(StateRegOutputF[108]) );
  XOR2_X1 F_StateRegOutput_Inst_LFInst_15_LFInst_4_U1 ( .A(StateRegOutput[61]), 
        .B(StateRegOutput[62]), .Z(StateRegOutputF[109]) );
  XOR2_X1 F_StateRegOutput_Inst_LFInst_15_LFInst_5_U1 ( .A(StateRegOutput[61]), 
        .B(StateRegOutput[63]), .Z(StateRegOutputF[110]) );
  XOR2_X1 F_StateRegOutput_Inst_LFInst_15_LFInst_6_U1 ( .A(StateRegOutput[62]), 
        .B(StateRegOutput[63]), .Z(StateRegOutputF[111]) );
  XOR2_X2 CipherErrorVecGen_XORInst_0_0_U1 ( .A(StateRegOutputF[0]), .B(
        Red_StateRegOutput[0]), .Z(CipherErrorVec[0]) );
  XOR2_X1 CipherErrorVecGen_XORInst_0_1_U1 ( .A(StateRegOutputF[1]), .B(
        Red_StateRegOutput[1]), .Z(CipherErrorVec[1]) );
  XOR2_X1 CipherErrorVecGen_XORInst_0_2_U1 ( .A(StateRegOutputF[2]), .B(
        Red_StateRegOutput[2]), .Z(CipherErrorVec[2]) );
  XOR2_X1 CipherErrorVecGen_XORInst_0_3_U2 ( .A(StateRegOutputF[3]), .B(
        Red_StateRegOutput[3]), .Z(CipherErrorVecGen_XORInst_0_3_n4) );
  BUF_X1 CipherErrorVecGen_XORInst_0_3_U1 ( .A(
        CipherErrorVecGen_XORInst_0_3_n4), .Z(CipherErrorVec[3]) );
  XOR2_X1 CipherErrorVecGen_XORInst_0_4_U1 ( .A(StateRegOutputF[4]), .B(
        Red_StateRegOutput[4]), .Z(CipherErrorVec[4]) );
  XOR2_X1 CipherErrorVecGen_XORInst_0_5_U1 ( .A(StateRegOutputF[5]), .B(
        Red_StateRegOutput[5]), .Z(CipherErrorVec[5]) );
  XOR2_X2 CipherErrorVecGen_XORInst_0_6_U1 ( .A(StateRegOutputF[6]), .B(
        Red_StateRegOutput[6]), .Z(CipherErrorVec[6]) );
  XOR2_X2 CipherErrorVecGen_XORInst_1_0_U1 ( .A(StateRegOutputF[7]), .B(
        Red_StateRegOutput[7]), .Z(CipherErrorVec[7]) );
  XOR2_X1 CipherErrorVecGen_XORInst_1_1_U1 ( .A(StateRegOutputF[8]), .B(
        Red_StateRegOutput[8]), .Z(CipherErrorVec[8]) );
  XOR2_X1 CipherErrorVecGen_XORInst_1_2_U1 ( .A(StateRegOutputF[9]), .B(
        Red_StateRegOutput[9]), .Z(CipherErrorVec[9]) );
  XOR2_X1 CipherErrorVecGen_XORInst_1_3_U2 ( .A(StateRegOutputF[10]), .B(
        Red_StateRegOutput[10]), .Z(CipherErrorVecGen_XORInst_1_3_n4) );
  BUF_X1 CipherErrorVecGen_XORInst_1_3_U1 ( .A(
        CipherErrorVecGen_XORInst_1_3_n4), .Z(CipherErrorVec[10]) );
  XOR2_X1 CipherErrorVecGen_XORInst_1_4_U1 ( .A(StateRegOutputF[11]), .B(
        Red_StateRegOutput[11]), .Z(CipherErrorVec[11]) );
  XOR2_X1 CipherErrorVecGen_XORInst_1_5_U1 ( .A(StateRegOutputF[12]), .B(
        Red_StateRegOutput[12]), .Z(CipherErrorVec[12]) );
  XOR2_X2 CipherErrorVecGen_XORInst_1_6_U1 ( .A(StateRegOutputF[13]), .B(
        Red_StateRegOutput[13]), .Z(CipherErrorVec[13]) );
  XOR2_X2 CipherErrorVecGen_XORInst_2_0_U1 ( .A(StateRegOutputF[14]), .B(
        Red_StateRegOutput[14]), .Z(CipherErrorVec[14]) );
  XOR2_X1 CipherErrorVecGen_XORInst_2_1_U1 ( .A(StateRegOutputF[15]), .B(
        Red_StateRegOutput[15]), .Z(CipherErrorVec[15]) );
  XOR2_X1 CipherErrorVecGen_XORInst_2_2_U1 ( .A(StateRegOutputF[16]), .B(
        Red_StateRegOutput[16]), .Z(CipherErrorVec[16]) );
  XOR2_X1 CipherErrorVecGen_XORInst_2_3_U2 ( .A(StateRegOutputF[17]), .B(
        Red_StateRegOutput[17]), .Z(CipherErrorVecGen_XORInst_2_3_n4) );
  BUF_X1 CipherErrorVecGen_XORInst_2_3_U1 ( .A(
        CipherErrorVecGen_XORInst_2_3_n4), .Z(CipherErrorVec[17]) );
  XOR2_X1 CipherErrorVecGen_XORInst_2_4_U1 ( .A(StateRegOutputF[18]), .B(
        Red_StateRegOutput[18]), .Z(CipherErrorVec[18]) );
  XOR2_X1 CipherErrorVecGen_XORInst_2_5_U1 ( .A(StateRegOutputF[19]), .B(
        Red_StateRegOutput[19]), .Z(CipherErrorVec[19]) );
  XOR2_X2 CipherErrorVecGen_XORInst_2_6_U1 ( .A(StateRegOutputF[20]), .B(
        Red_StateRegOutput[20]), .Z(CipherErrorVec[20]) );
  XOR2_X2 CipherErrorVecGen_XORInst_3_0_U1 ( .A(StateRegOutputF[21]), .B(
        Red_StateRegOutput[21]), .Z(CipherErrorVec[21]) );
  XOR2_X1 CipherErrorVecGen_XORInst_3_1_U1 ( .A(StateRegOutputF[22]), .B(
        Red_StateRegOutput[22]), .Z(CipherErrorVec[22]) );
  XOR2_X1 CipherErrorVecGen_XORInst_3_2_U1 ( .A(StateRegOutputF[23]), .B(
        Red_StateRegOutput[23]), .Z(CipherErrorVec[23]) );
  XOR2_X1 CipherErrorVecGen_XORInst_3_3_U2 ( .A(StateRegOutputF[24]), .B(
        Red_StateRegOutput[24]), .Z(CipherErrorVecGen_XORInst_3_3_n4) );
  BUF_X1 CipherErrorVecGen_XORInst_3_3_U1 ( .A(
        CipherErrorVecGen_XORInst_3_3_n4), .Z(CipherErrorVec[24]) );
  XOR2_X1 CipherErrorVecGen_XORInst_3_4_U1 ( .A(StateRegOutputF[25]), .B(
        Red_StateRegOutput[25]), .Z(CipherErrorVec[25]) );
  XOR2_X1 CipherErrorVecGen_XORInst_3_5_U1 ( .A(StateRegOutputF[26]), .B(
        Red_StateRegOutput[26]), .Z(CipherErrorVec[26]) );
  XOR2_X2 CipherErrorVecGen_XORInst_3_6_U1 ( .A(StateRegOutputF[27]), .B(
        Red_StateRegOutput[27]), .Z(CipherErrorVec[27]) );
  XOR2_X2 CipherErrorVecGen_XORInst_4_0_U1 ( .A(StateRegOutputF[28]), .B(
        Red_StateRegOutput[28]), .Z(CipherErrorVec[28]) );
  XOR2_X1 CipherErrorVecGen_XORInst_4_1_U1 ( .A(StateRegOutputF[29]), .B(
        Red_StateRegOutput[29]), .Z(CipherErrorVec[29]) );
  XOR2_X1 CipherErrorVecGen_XORInst_4_2_U1 ( .A(StateRegOutputF[30]), .B(
        Red_StateRegOutput[30]), .Z(CipherErrorVec[30]) );
  XOR2_X1 CipherErrorVecGen_XORInst_4_3_U2 ( .A(StateRegOutputF[31]), .B(
        Red_StateRegOutput[31]), .Z(CipherErrorVecGen_XORInst_4_3_n4) );
  BUF_X1 CipherErrorVecGen_XORInst_4_3_U1 ( .A(
        CipherErrorVecGen_XORInst_4_3_n4), .Z(CipherErrorVec[31]) );
  XOR2_X1 CipherErrorVecGen_XORInst_4_4_U1 ( .A(StateRegOutputF[32]), .B(
        Red_StateRegOutput[32]), .Z(CipherErrorVec[32]) );
  XOR2_X1 CipherErrorVecGen_XORInst_4_5_U1 ( .A(StateRegOutputF[33]), .B(
        Red_StateRegOutput[33]), .Z(CipherErrorVec[33]) );
  XOR2_X2 CipherErrorVecGen_XORInst_4_6_U1 ( .A(StateRegOutputF[34]), .B(
        Red_StateRegOutput[34]), .Z(CipherErrorVec[34]) );
  XOR2_X2 CipherErrorVecGen_XORInst_5_0_U1 ( .A(StateRegOutputF[35]), .B(
        Red_StateRegOutput[35]), .Z(CipherErrorVec[35]) );
  XOR2_X1 CipherErrorVecGen_XORInst_5_1_U1 ( .A(StateRegOutputF[36]), .B(
        Red_StateRegOutput[36]), .Z(CipherErrorVec[36]) );
  XOR2_X1 CipherErrorVecGen_XORInst_5_2_U1 ( .A(StateRegOutputF[37]), .B(
        Red_StateRegOutput[37]), .Z(CipherErrorVec[37]) );
  XOR2_X1 CipherErrorVecGen_XORInst_5_3_U2 ( .A(StateRegOutputF[38]), .B(
        Red_StateRegOutput[38]), .Z(CipherErrorVecGen_XORInst_5_3_n4) );
  BUF_X1 CipherErrorVecGen_XORInst_5_3_U1 ( .A(
        CipherErrorVecGen_XORInst_5_3_n4), .Z(CipherErrorVec[38]) );
  XOR2_X1 CipherErrorVecGen_XORInst_5_4_U1 ( .A(StateRegOutputF[39]), .B(
        Red_StateRegOutput[39]), .Z(CipherErrorVec[39]) );
  XOR2_X1 CipherErrorVecGen_XORInst_5_5_U1 ( .A(StateRegOutputF[40]), .B(
        Red_StateRegOutput[40]), .Z(CipherErrorVec[40]) );
  XOR2_X2 CipherErrorVecGen_XORInst_5_6_U1 ( .A(StateRegOutputF[41]), .B(
        Red_StateRegOutput[41]), .Z(CipherErrorVec[41]) );
  XOR2_X2 CipherErrorVecGen_XORInst_6_0_U1 ( .A(StateRegOutputF[42]), .B(
        Red_StateRegOutput[42]), .Z(CipherErrorVec[42]) );
  XOR2_X1 CipherErrorVecGen_XORInst_6_1_U1 ( .A(StateRegOutputF[43]), .B(
        Red_StateRegOutput[43]), .Z(CipherErrorVec[43]) );
  XOR2_X1 CipherErrorVecGen_XORInst_6_2_U1 ( .A(StateRegOutputF[44]), .B(
        Red_StateRegOutput[44]), .Z(CipherErrorVec[44]) );
  XOR2_X1 CipherErrorVecGen_XORInst_6_3_U2 ( .A(StateRegOutputF[45]), .B(
        Red_StateRegOutput[45]), .Z(CipherErrorVecGen_XORInst_6_3_n4) );
  BUF_X1 CipherErrorVecGen_XORInst_6_3_U1 ( .A(
        CipherErrorVecGen_XORInst_6_3_n4), .Z(CipherErrorVec[45]) );
  XOR2_X1 CipherErrorVecGen_XORInst_6_4_U1 ( .A(StateRegOutputF[46]), .B(
        Red_StateRegOutput[46]), .Z(CipherErrorVec[46]) );
  XOR2_X1 CipherErrorVecGen_XORInst_6_5_U1 ( .A(StateRegOutputF[47]), .B(
        Red_StateRegOutput[47]), .Z(CipherErrorVec[47]) );
  XOR2_X2 CipherErrorVecGen_XORInst_6_6_U1 ( .A(StateRegOutputF[48]), .B(
        Red_StateRegOutput[48]), .Z(CipherErrorVec[48]) );
  XOR2_X2 CipherErrorVecGen_XORInst_7_0_U1 ( .A(StateRegOutputF[49]), .B(
        Red_StateRegOutput[49]), .Z(CipherErrorVec[49]) );
  XOR2_X1 CipherErrorVecGen_XORInst_7_1_U1 ( .A(StateRegOutputF[50]), .B(
        Red_StateRegOutput[50]), .Z(CipherErrorVec[50]) );
  XOR2_X1 CipherErrorVecGen_XORInst_7_2_U1 ( .A(StateRegOutputF[51]), .B(
        Red_StateRegOutput[51]), .Z(CipherErrorVec[51]) );
  XOR2_X1 CipherErrorVecGen_XORInst_7_3_U2 ( .A(StateRegOutputF[52]), .B(
        Red_StateRegOutput[52]), .Z(CipherErrorVecGen_XORInst_7_3_n4) );
  BUF_X1 CipherErrorVecGen_XORInst_7_3_U1 ( .A(
        CipherErrorVecGen_XORInst_7_3_n4), .Z(CipherErrorVec[52]) );
  XOR2_X1 CipherErrorVecGen_XORInst_7_4_U1 ( .A(StateRegOutputF[53]), .B(
        Red_StateRegOutput[53]), .Z(CipherErrorVec[53]) );
  XOR2_X1 CipherErrorVecGen_XORInst_7_5_U1 ( .A(StateRegOutputF[54]), .B(
        Red_StateRegOutput[54]), .Z(CipherErrorVec[54]) );
  XOR2_X2 CipherErrorVecGen_XORInst_7_6_U1 ( .A(StateRegOutputF[55]), .B(
        Red_StateRegOutput[55]), .Z(CipherErrorVec[55]) );
  XOR2_X2 CipherErrorVecGen_XORInst_8_0_U1 ( .A(StateRegOutputF[56]), .B(
        Red_StateRegOutput[56]), .Z(CipherErrorVec[56]) );
  XOR2_X1 CipherErrorVecGen_XORInst_8_1_U1 ( .A(StateRegOutputF[57]), .B(
        Red_StateRegOutput[57]), .Z(CipherErrorVec[57]) );
  XOR2_X1 CipherErrorVecGen_XORInst_8_2_U1 ( .A(StateRegOutputF[58]), .B(
        Red_StateRegOutput[58]), .Z(CipherErrorVec[58]) );
  XOR2_X1 CipherErrorVecGen_XORInst_8_3_U2 ( .A(StateRegOutputF[59]), .B(
        Red_StateRegOutput[59]), .Z(CipherErrorVecGen_XORInst_8_3_n4) );
  BUF_X1 CipherErrorVecGen_XORInst_8_3_U1 ( .A(
        CipherErrorVecGen_XORInst_8_3_n4), .Z(CipherErrorVec[59]) );
  XOR2_X1 CipherErrorVecGen_XORInst_8_4_U1 ( .A(StateRegOutputF[60]), .B(
        Red_StateRegOutput[60]), .Z(CipherErrorVec[60]) );
  XOR2_X1 CipherErrorVecGen_XORInst_8_5_U1 ( .A(StateRegOutputF[61]), .B(
        Red_StateRegOutput[61]), .Z(CipherErrorVec[61]) );
  XOR2_X2 CipherErrorVecGen_XORInst_8_6_U1 ( .A(StateRegOutputF[62]), .B(
        Red_StateRegOutput[62]), .Z(CipherErrorVec[62]) );
  XOR2_X2 CipherErrorVecGen_XORInst_9_0_U1 ( .A(StateRegOutputF[63]), .B(
        Red_StateRegOutput[63]), .Z(CipherErrorVec[63]) );
  XOR2_X1 CipherErrorVecGen_XORInst_9_1_U1 ( .A(StateRegOutputF[64]), .B(
        Red_StateRegOutput[64]), .Z(CipherErrorVec[64]) );
  XOR2_X1 CipherErrorVecGen_XORInst_9_2_U1 ( .A(StateRegOutputF[65]), .B(
        Red_StateRegOutput[65]), .Z(CipherErrorVec[65]) );
  XOR2_X1 CipherErrorVecGen_XORInst_9_3_U2 ( .A(StateRegOutputF[66]), .B(
        Red_StateRegOutput[66]), .Z(CipherErrorVecGen_XORInst_9_3_n4) );
  BUF_X1 CipherErrorVecGen_XORInst_9_3_U1 ( .A(
        CipherErrorVecGen_XORInst_9_3_n4), .Z(CipherErrorVec[66]) );
  XOR2_X1 CipherErrorVecGen_XORInst_9_4_U1 ( .A(StateRegOutputF[67]), .B(
        Red_StateRegOutput[67]), .Z(CipherErrorVec[67]) );
  XOR2_X1 CipherErrorVecGen_XORInst_9_5_U1 ( .A(StateRegOutputF[68]), .B(
        Red_StateRegOutput[68]), .Z(CipherErrorVec[68]) );
  XOR2_X2 CipherErrorVecGen_XORInst_9_6_U1 ( .A(StateRegOutputF[69]), .B(
        Red_StateRegOutput[69]), .Z(CipherErrorVec[69]) );
  XOR2_X2 CipherErrorVecGen_XORInst_10_0_U1 ( .A(StateRegOutputF[70]), .B(
        Red_StateRegOutput[70]), .Z(CipherErrorVec[70]) );
  XOR2_X1 CipherErrorVecGen_XORInst_10_1_U1 ( .A(StateRegOutputF[71]), .B(
        Red_StateRegOutput[71]), .Z(CipherErrorVec[71]) );
  XOR2_X1 CipherErrorVecGen_XORInst_10_2_U1 ( .A(StateRegOutputF[72]), .B(
        Red_StateRegOutput[72]), .Z(CipherErrorVec[72]) );
  XOR2_X1 CipherErrorVecGen_XORInst_10_3_U2 ( .A(StateRegOutputF[73]), .B(
        Red_StateRegOutput[73]), .Z(CipherErrorVecGen_XORInst_10_3_n4) );
  BUF_X1 CipherErrorVecGen_XORInst_10_3_U1 ( .A(
        CipherErrorVecGen_XORInst_10_3_n4), .Z(CipherErrorVec[73]) );
  XOR2_X1 CipherErrorVecGen_XORInst_10_4_U1 ( .A(StateRegOutputF[74]), .B(
        Red_StateRegOutput[74]), .Z(CipherErrorVec[74]) );
  XOR2_X1 CipherErrorVecGen_XORInst_10_5_U1 ( .A(StateRegOutputF[75]), .B(
        Red_StateRegOutput[75]), .Z(CipherErrorVec[75]) );
  XOR2_X2 CipherErrorVecGen_XORInst_10_6_U1 ( .A(StateRegOutputF[76]), .B(
        Red_StateRegOutput[76]), .Z(CipherErrorVec[76]) );
  XOR2_X2 CipherErrorVecGen_XORInst_11_0_U1 ( .A(StateRegOutputF[77]), .B(
        Red_StateRegOutput[77]), .Z(CipherErrorVec[77]) );
  XOR2_X1 CipherErrorVecGen_XORInst_11_1_U1 ( .A(StateRegOutputF[78]), .B(
        Red_StateRegOutput[78]), .Z(CipherErrorVec[78]) );
  XOR2_X1 CipherErrorVecGen_XORInst_11_2_U1 ( .A(StateRegOutputF[79]), .B(
        Red_StateRegOutput[79]), .Z(CipherErrorVec[79]) );
  XOR2_X1 CipherErrorVecGen_XORInst_11_3_U2 ( .A(StateRegOutputF[80]), .B(
        Red_StateRegOutput[80]), .Z(CipherErrorVecGen_XORInst_11_3_n4) );
  BUF_X1 CipherErrorVecGen_XORInst_11_3_U1 ( .A(
        CipherErrorVecGen_XORInst_11_3_n4), .Z(CipherErrorVec[80]) );
  XOR2_X1 CipherErrorVecGen_XORInst_11_4_U1 ( .A(StateRegOutputF[81]), .B(
        Red_StateRegOutput[81]), .Z(CipherErrorVec[81]) );
  XOR2_X1 CipherErrorVecGen_XORInst_11_5_U1 ( .A(StateRegOutputF[82]), .B(
        Red_StateRegOutput[82]), .Z(CipherErrorVec[82]) );
  XOR2_X2 CipherErrorVecGen_XORInst_11_6_U1 ( .A(StateRegOutputF[83]), .B(
        Red_StateRegOutput[83]), .Z(CipherErrorVec[83]) );
  XOR2_X2 CipherErrorVecGen_XORInst_12_0_U1 ( .A(StateRegOutputF[84]), .B(
        Red_StateRegOutput[84]), .Z(CipherErrorVec[84]) );
  XOR2_X1 CipherErrorVecGen_XORInst_12_1_U1 ( .A(StateRegOutputF[85]), .B(
        Red_StateRegOutput[85]), .Z(CipherErrorVec[85]) );
  XOR2_X1 CipherErrorVecGen_XORInst_12_2_U1 ( .A(StateRegOutputF[86]), .B(
        Red_StateRegOutput[86]), .Z(CipherErrorVec[86]) );
  XOR2_X1 CipherErrorVecGen_XORInst_12_3_U2 ( .A(StateRegOutputF[87]), .B(
        Red_StateRegOutput[87]), .Z(CipherErrorVecGen_XORInst_12_3_n4) );
  BUF_X1 CipherErrorVecGen_XORInst_12_3_U1 ( .A(
        CipherErrorVecGen_XORInst_12_3_n4), .Z(CipherErrorVec[87]) );
  XOR2_X1 CipherErrorVecGen_XORInst_12_4_U1 ( .A(StateRegOutputF[88]), .B(
        Red_StateRegOutput[88]), .Z(CipherErrorVec[88]) );
  XOR2_X1 CipherErrorVecGen_XORInst_12_5_U1 ( .A(StateRegOutputF[89]), .B(
        Red_StateRegOutput[89]), .Z(CipherErrorVec[89]) );
  XOR2_X2 CipherErrorVecGen_XORInst_12_6_U1 ( .A(StateRegOutputF[90]), .B(
        Red_StateRegOutput[90]), .Z(CipherErrorVec[90]) );
  XOR2_X2 CipherErrorVecGen_XORInst_13_0_U1 ( .A(StateRegOutputF[91]), .B(
        Red_StateRegOutput[91]), .Z(CipherErrorVec[91]) );
  XOR2_X1 CipherErrorVecGen_XORInst_13_1_U1 ( .A(StateRegOutputF[92]), .B(
        Red_StateRegOutput[92]), .Z(CipherErrorVec[92]) );
  XOR2_X1 CipherErrorVecGen_XORInst_13_2_U1 ( .A(StateRegOutputF[93]), .B(
        Red_StateRegOutput[93]), .Z(CipherErrorVec[93]) );
  XOR2_X1 CipherErrorVecGen_XORInst_13_3_U2 ( .A(StateRegOutputF[94]), .B(
        Red_StateRegOutput[94]), .Z(CipherErrorVecGen_XORInst_13_3_n4) );
  BUF_X1 CipherErrorVecGen_XORInst_13_3_U1 ( .A(
        CipherErrorVecGen_XORInst_13_3_n4), .Z(CipherErrorVec[94]) );
  XOR2_X1 CipherErrorVecGen_XORInst_13_4_U1 ( .A(StateRegOutputF[95]), .B(
        Red_StateRegOutput[95]), .Z(CipherErrorVec[95]) );
  XOR2_X1 CipherErrorVecGen_XORInst_13_5_U1 ( .A(StateRegOutputF[96]), .B(
        Red_StateRegOutput[96]), .Z(CipherErrorVec[96]) );
  XOR2_X2 CipherErrorVecGen_XORInst_13_6_U1 ( .A(StateRegOutputF[97]), .B(
        Red_StateRegOutput[97]), .Z(CipherErrorVec[97]) );
  XOR2_X2 CipherErrorVecGen_XORInst_14_0_U1 ( .A(StateRegOutputF[98]), .B(
        Red_StateRegOutput[98]), .Z(CipherErrorVec[98]) );
  XOR2_X1 CipherErrorVecGen_XORInst_14_1_U1 ( .A(StateRegOutputF[99]), .B(
        Red_StateRegOutput[99]), .Z(CipherErrorVec[99]) );
  XOR2_X1 CipherErrorVecGen_XORInst_14_2_U1 ( .A(StateRegOutputF[100]), .B(
        Red_StateRegOutput[100]), .Z(CipherErrorVec[100]) );
  XOR2_X1 CipherErrorVecGen_XORInst_14_3_U2 ( .A(StateRegOutputF[101]), .B(
        Red_StateRegOutput[101]), .Z(CipherErrorVecGen_XORInst_14_3_n4) );
  BUF_X1 CipherErrorVecGen_XORInst_14_3_U1 ( .A(
        CipherErrorVecGen_XORInst_14_3_n4), .Z(CipherErrorVec[101]) );
  XOR2_X1 CipherErrorVecGen_XORInst_14_4_U1 ( .A(StateRegOutputF[102]), .B(
        Red_StateRegOutput[102]), .Z(CipherErrorVec[102]) );
  XOR2_X1 CipherErrorVecGen_XORInst_14_5_U1 ( .A(StateRegOutputF[103]), .B(
        Red_StateRegOutput[103]), .Z(CipherErrorVec[103]) );
  XOR2_X2 CipherErrorVecGen_XORInst_14_6_U1 ( .A(StateRegOutputF[104]), .B(
        Red_StateRegOutput[104]), .Z(CipherErrorVec[104]) );
  XOR2_X2 CipherErrorVecGen_XORInst_15_0_U1 ( .A(StateRegOutputF[105]), .B(
        Red_StateRegOutput[105]), .Z(CipherErrorVec[105]) );
  XOR2_X1 CipherErrorVecGen_XORInst_15_1_U1 ( .A(StateRegOutputF[106]), .B(
        Red_StateRegOutput[106]), .Z(CipherErrorVec[106]) );
  XOR2_X1 CipherErrorVecGen_XORInst_15_2_U1 ( .A(StateRegOutputF[107]), .B(
        Red_StateRegOutput[107]), .Z(CipherErrorVec[107]) );
  XOR2_X1 CipherErrorVecGen_XORInst_15_3_U2 ( .A(StateRegOutputF[108]), .B(
        Red_StateRegOutput[108]), .Z(CipherErrorVecGen_XORInst_15_3_n4) );
  BUF_X1 CipherErrorVecGen_XORInst_15_3_U1 ( .A(
        CipherErrorVecGen_XORInst_15_3_n4), .Z(CipherErrorVec[108]) );
  XOR2_X1 CipherErrorVecGen_XORInst_15_4_U1 ( .A(StateRegOutputF[109]), .B(
        Red_StateRegOutput[109]), .Z(CipherErrorVec[109]) );
  XOR2_X1 CipherErrorVecGen_XORInst_15_5_U1 ( .A(StateRegOutputF[110]), .B(
        Red_StateRegOutput[110]), .Z(CipherErrorVec[110]) );
  XOR2_X2 CipherErrorVecGen_XORInst_15_6_U1 ( .A(StateRegOutputF[111]), .B(
        Red_StateRegOutput[111]), .Z(CipherErrorVec[111]) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_0_U47 ( .B1(OutputRegIn[2]), .B2(
        OutputRegIn[3]), .A(SD1_SB_inst_SD1_SB_bit_inst_0_n131), .ZN(
        Feedback[60]) );
  AOI221_X1 SD1_SB_inst_SD1_SB_bit_inst_0_U46 ( .B1(OutputRegIn[2]), .B2(
        OutputRegIn[0]), .C1(OutputRegIn[3]), .C2(OutputRegIn[0]), .A(
        OutputRegIn[1]), .ZN(SD1_SB_inst_SD1_SB_bit_inst_0_n131) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_0_U45 ( .A(StateRegOutput[3]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_0_n127), .ZN(OutputRegIn[3]) );
  AOI211_X1 SD1_SB_inst_SD1_SB_bit_inst_0_U44 ( .C1(CipherErrorVec[6]), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_0_n126), .A(
        SD1_SB_inst_SD1_SB_bit_inst_0_n125), .B(
        SD1_SB_inst_SD1_SB_bit_inst_0_n124), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_0_n127) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_0_U43 ( .A1(CipherErrorVec[0]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_0_n101), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_0_n123), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_0_n124) );
  AOI222_X1 SD1_SB_inst_SD1_SB_bit_inst_0_U42 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_0_n108), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_0_n104), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_0_n108), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_0_n122), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_0_n104), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_0_n121), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_0_n126) );
  OAI221_X1 SD1_SB_inst_SD1_SB_bit_inst_0_U41 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_0_n120), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_0_n100), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_0_n120), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_0_n102), .A(
        SD1_SB_inst_SD1_SB_bit_inst_0_n106), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_0_n121) );
  OAI211_X1 SD1_SB_inst_SD1_SB_bit_inst_0_U40 ( .C1(
        SD1_SB_inst_SD1_SB_bit_inst_0_n105), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_0_n100), .A(
        SD1_SB_inst_SD1_SB_bit_inst_0_n119), .B(
        SD1_SB_inst_SD1_SB_bit_inst_0_n102), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_0_n122) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_0_U39 ( .A(StateRegOutput[2]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_0_n118), .ZN(OutputRegIn[2]) );
  AOI211_X1 SD1_SB_inst_SD1_SB_bit_inst_0_U38 ( .C1(CipherErrorVec[6]), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_0_n117), .A(
        SD1_SB_inst_SD1_SB_bit_inst_0_n125), .B(
        SD1_SB_inst_SD1_SB_bit_inst_0_n116), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_0_n118) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_0_U37 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_0_n128), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_0_n96), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_0_n116) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_0_U36 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_0_n105), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_0_n120), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_0_n128) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_0_U35 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_0_n102), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_0_n123), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_0_n119), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_0_n125) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_0_U34 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_0_n105), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_0_n100), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_0_n119) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_0_U33 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_0_n107), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_0_n103), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_0_n123) );
  OAI22_X1 SD1_SB_inst_SD1_SB_bit_inst_0_U32 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_0_n107), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_0_n115), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_0_n114), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_0_n102), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_0_n117) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_0_U31 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_0_n100), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_0_n104), .A(
        SD1_SB_inst_SD1_SB_bit_inst_0_n105), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_0_n114) );
  AOI22_X1 SD1_SB_inst_SD1_SB_bit_inst_0_U30 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_0_n105), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_0_n100), .B1(CipherErrorVec[0]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_0_n113), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_0_n115) );
  OAI21_X1 SD1_SB_inst_SD1_SB_bit_inst_0_U29 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_0_n103), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_0_n106), .A(
        SD1_SB_inst_SD1_SB_bit_inst_0_n112), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_0_n113) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_0_U28 ( .A(StateRegOutput[0]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_0_n111), .ZN(OutputRegIn[0]) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_0_U27 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_0_n110), .B2(CipherErrorVec[2]), .A(
        SD1_SB_inst_SD1_SB_bit_inst_0_n109), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_0_n111) );
  AOI221_X1 SD1_SB_inst_SD1_SB_bit_inst_0_U26 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_0_n107), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_0_n112), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_0_n108), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_0_n129), .A(
        SD1_SB_inst_SD1_SB_bit_inst_0_n104), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_0_n109) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_0_U25 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_0_n120), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_0_n112) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_0_U24 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_0_n100), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_0_n102), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_0_n120) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_0_U23 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_0_n130), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_0_n105), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_0_n110) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_0_U22 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_0_n108), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_0_n107) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_0_U21 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_0_n106), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_0_n105) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_0_U20 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_0_n104), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_0_n103) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_0_U19 ( .A(CipherErrorVec[2]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_0_n102) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_0_U18 ( .A(CipherErrorVec[1]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_0_n101) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_0_U17 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_0_n101), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_0_n100) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_0_U16 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_0_n99), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_0_n130) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_0_U15 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_0_n97), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_0_n129) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_0_U14 ( .A(CipherErrorVec[0]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_0_n96) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_0_U13 ( .A(CipherErrorVec[5]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_0_n108) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_0_U12 ( .A(CipherErrorVec[4]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_0_n106) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_0_U11 ( .A(CipherErrorVec[3]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_0_n104) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_0_U10 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_0_n100), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_0_n107), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_0_n98) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_0_U9 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_0_n98), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_0_n104), .A(
        SD1_SB_inst_SD1_SB_bit_inst_0_n96), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_0_n99) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_0_U8 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_0_n105), .A2(CipherErrorVec[2]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_0_n95) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_0_U7 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_0_n95), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_0_n96), .A(
        SD1_SB_inst_SD1_SB_bit_inst_0_n101), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_0_n97) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_0_U6 ( .A(StateRegOutput[1]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_0_n94), .ZN(OutputRegIn[1]) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_0_U5 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_0_n107), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_0_n92), .A(
        SD1_SB_inst_SD1_SB_bit_inst_0_n93), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_0_n94) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_0_U4 ( .A1(CipherErrorVec[2]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_0_n130), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_0_n106), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_0_n93) );
  OAI22_X1 SD1_SB_inst_SD1_SB_bit_inst_0_U3 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_0_n103), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_0_n129), .B1(CipherErrorVec[6]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_0_n128), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_0_n92) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_1_U37 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_1_n110), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_1_n109), .A(
        SD1_SB_inst_SD1_SB_bit_inst_1_n108), .ZN(Feedback[61]) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_1_U36 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_1_n107), .B2(StateRegOutput[0]), .A(
        SD1_SB_inst_SD1_SB_bit_inst_1_n106), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_1_n108) );
  OAI22_X1 SD1_SB_inst_SD1_SB_bit_inst_1_U35 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_1_n109), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_1_n110), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_1_n107), .B2(StateRegOutput[0]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_1_n106) );
  AOI22_X1 SD1_SB_inst_SD1_SB_bit_inst_1_U34 ( .A1(CipherErrorVec[0]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_1_n105), .B1(CipherErrorVec[3]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_1_n104), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_1_n107) );
  OAI21_X1 SD1_SB_inst_SD1_SB_bit_inst_1_U33 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_1_n103), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_1_n102), .A(
        SD1_SB_inst_SD1_SB_bit_inst_1_n101), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_1_n104) );
  NAND3_X1 SD1_SB_inst_SD1_SB_bit_inst_1_U32 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_1_n79), .A2(CipherErrorVec[5]), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_1_n78), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_1_n101) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_1_U31 ( .A1(CipherErrorVec[0]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_1_n79), .A3(CipherErrorVec[4]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_1_n103) );
  AOI211_X1 SD1_SB_inst_SD1_SB_bit_inst_1_U30 ( .C1(
        SD1_SB_inst_SD1_SB_bit_inst_1_n100), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_1_n78), .A(CipherErrorVec[4]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_1_n80), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_1_n105) );
  XOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_1_U29 ( .A(StateRegOutput[2]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_1_n99), .Z(
        SD1_SB_inst_SD1_SB_bit_inst_1_n109) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_1_U28 ( .B1(CipherErrorVec[6]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_1_n98), .A(
        SD1_SB_inst_SD1_SB_bit_inst_1_n97), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_1_n99) );
  AOI221_X1 SD1_SB_inst_SD1_SB_bit_inst_1_U27 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_1_n77), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_1_n96), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_1_n78), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_1_n95), .A(
        SD1_SB_inst_SD1_SB_bit_inst_1_n94), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_1_n97) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_1_U26 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_1_n93), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_1_n94) );
  OAI22_X1 SD1_SB_inst_SD1_SB_bit_inst_1_U25 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_1_n92), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_1_n80), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_1_n91), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_1_n82), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_1_n98) );
  AOI211_X1 SD1_SB_inst_SD1_SB_bit_inst_1_U24 ( .C1(CipherErrorVec[0]), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_1_n100), .A(
        SD1_SB_inst_SD1_SB_bit_inst_1_n79), .B(
        SD1_SB_inst_SD1_SB_bit_inst_1_n90), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_1_n91) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_1_U23 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_1_n102), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_1_n90) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_1_U22 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_1_n77), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_1_n83), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_1_n102) );
  AOI22_X1 SD1_SB_inst_SD1_SB_bit_inst_1_U21 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_1_n77), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_1_n81), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_1_n89), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_1_n83), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_1_n92) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_1_U20 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_1_n77), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_1_n95), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_1_n89) );
  XOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_1_U19 ( .A(StateRegOutput[3]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_1_n88), .Z(
        SD1_SB_inst_SD1_SB_bit_inst_1_n110) );
  OAI21_X1 SD1_SB_inst_SD1_SB_bit_inst_1_U18 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_1_n87), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_1_n96), .A(
        SD1_SB_inst_SD1_SB_bit_inst_1_n86), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_1_n88) );
  OAI221_X1 SD1_SB_inst_SD1_SB_bit_inst_1_U17 ( .B1(CipherErrorVec[4]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_1_n85), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_1_n82), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_1_n84), .A(CipherErrorVec[6]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_1_n86) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_1_U16 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_1_n77), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_1_n79), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_1_n81), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_1_n84) );
  OAI33_X1 SD1_SB_inst_SD1_SB_bit_inst_1_U15 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_1_n79), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_1_n100), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_1_n78), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_1_n80), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_1_n83), .B3(
        SD1_SB_inst_SD1_SB_bit_inst_1_n77), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_1_n85) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_1_U14 ( .A1(CipherErrorVec[3]), .A2(
        CipherErrorVec[5]), .ZN(SD1_SB_inst_SD1_SB_bit_inst_1_n100) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_1_U13 ( .A1(CipherErrorVec[3]), .A2(
        CipherErrorVec[5]), .ZN(SD1_SB_inst_SD1_SB_bit_inst_1_n96) );
  AOI221_X1 SD1_SB_inst_SD1_SB_bit_inst_1_U12 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_1_n93), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_1_n77), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_1_n95), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_1_n77), .A(CipherErrorVec[6]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_1_n87) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_1_U11 ( .A(CipherErrorVec[0]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_1_n95) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_1_U10 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_1_n80), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_1_n82), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_1_n93) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_1_U9 ( .A(CipherErrorVec[3]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_1_n81) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_1_U8 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_1_n80), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_1_n79) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_1_U7 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_1_n78), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_1_n77) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_1_U6 ( .A(CipherErrorVec[4]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_1_n82) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_1_U5 ( .A(CipherErrorVec[5]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_1_n83) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_1_U4 ( .A(CipherErrorVec[2]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_1_n80) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_1_U3 ( .A(CipherErrorVec[1]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_1_n78) );
  OAI22_X1 SD1_SB_inst_SD1_SB_bit_inst_2_U45 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_2_n138), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_2_n137), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_2_n136), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_2_n135), .ZN(Feedback[62]) );
  XOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_2_U44 ( .A(StateRegOutput[1]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_2_n134), .Z(
        SD1_SB_inst_SD1_SB_bit_inst_2_n137) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_2_U43 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_2_n103), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_2_n133), .A(
        SD1_SB_inst_SD1_SB_bit_inst_2_n132), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_2_n134) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_2_U42 ( .A1(CipherErrorVec[3]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_2_n131), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_2_n130), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_2_n132) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_2_U41 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_2_n105), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_2_n99), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_2_n130) );
  OAI22_X1 SD1_SB_inst_SD1_SB_bit_inst_2_U40 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_2_n101), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_2_n129), .B1(CipherErrorVec[6]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_2_n128), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_2_n133) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_2_U39 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_2_n135), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_2_n136), .A(
        SD1_SB_inst_SD1_SB_bit_inst_2_n127), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_2_n138) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_2_U38 ( .A(StateRegOutput[2]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_2_n126), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_2_n127) );
  AOI211_X1 SD1_SB_inst_SD1_SB_bit_inst_2_U37 ( .C1(
        SD1_SB_inst_SD1_SB_bit_inst_2_n101), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_2_n125), .A(
        SD1_SB_inst_SD1_SB_bit_inst_2_n124), .B(
        SD1_SB_inst_SD1_SB_bit_inst_2_n123), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_2_n126) );
  AOI211_X1 SD1_SB_inst_SD1_SB_bit_inst_2_U36 ( .C1(
        SD1_SB_inst_SD1_SB_bit_inst_2_n122), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_2_n102), .A(
        SD1_SB_inst_SD1_SB_bit_inst_2_n121), .B(
        SD1_SB_inst_SD1_SB_bit_inst_2_n104), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_2_n123) );
  AOI22_X1 SD1_SB_inst_SD1_SB_bit_inst_2_U35 ( .A1(CipherErrorVec[0]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_2_n120), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_2_n99), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_2_n106), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_2_n122) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_2_U34 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_2_n102), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_2_n104), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_2_n119), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_2_n124) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_2_U33 ( .A(CipherErrorVec[6]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_2_n121) );
  OAI221_X1 SD1_SB_inst_SD1_SB_bit_inst_2_U32 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_2_n103), .B2(CipherErrorVec[6]), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_2_n103), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_2_n106), .A(CipherErrorVec[0]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_2_n118) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_2_U31 ( .A(StateRegOutput[0]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_2_n117), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_2_n136) );
  AOI22_X1 SD1_SB_inst_SD1_SB_bit_inst_2_U30 ( .A1(CipherErrorVec[3]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_2_n116), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_2_n101), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_2_n115), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_2_n117) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_2_U29 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_2_n103), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_2_n129), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_2_n115) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_2_U28 ( .A1(CipherErrorVec[0]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_2_n114), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_2_n129) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_2_U27 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_2_n120), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_2_n100), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_2_n114) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_2_U26 ( .A1(CipherErrorVec[3]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_2_n105), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_2_n120) );
  OAI21_X1 SD1_SB_inst_SD1_SB_bit_inst_2_U25 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_2_n131), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_2_n113), .A(
        SD1_SB_inst_SD1_SB_bit_inst_2_n128), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_2_n116) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_2_U24 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_2_n99), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_2_n106), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_2_n113) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_2_U23 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_2_n101), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_2_n103), .A3(CipherErrorVec[0]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_2_n131) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_2_U22 ( .A(StateRegOutput[3]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_2_n112), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_2_n135) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_2_U21 ( .B1(CipherErrorVec[6]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_2_n111), .A(
        SD1_SB_inst_SD1_SB_bit_inst_2_n110), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_2_n112) );
  AOI221_X1 SD1_SB_inst_SD1_SB_bit_inst_2_U20 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_2_n104), .B2(CipherErrorVec[0]), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_2_n102), .C2(CipherErrorVec[0]), .A(
        SD1_SB_inst_SD1_SB_bit_inst_2_n119), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_2_n110) );
  NAND3_X1 SD1_SB_inst_SD1_SB_bit_inst_2_U19 ( .A1(CipherErrorVec[3]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_2_n105), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_2_n99), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_2_n119) );
  OAI221_X1 SD1_SB_inst_SD1_SB_bit_inst_2_U18 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_2_n103), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_2_n128), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_2_n103), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_2_n109), .A(
        SD1_SB_inst_SD1_SB_bit_inst_2_n108), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_2_n111) );
  OAI21_X1 SD1_SB_inst_SD1_SB_bit_inst_2_U17 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_2_n105), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_2_n107), .A(CipherErrorVec[3]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_2_n108) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_2_U16 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_2_n101), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_2_n99), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_2_n104), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_2_n107) );
  OAI211_X1 SD1_SB_inst_SD1_SB_bit_inst_2_U15 ( .C1(CipherErrorVec[3]), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_2_n105), .A(
        SD1_SB_inst_SD1_SB_bit_inst_2_n99), .B(
        SD1_SB_inst_SD1_SB_bit_inst_2_n102), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_2_n109) );
  NAND3_X1 SD1_SB_inst_SD1_SB_bit_inst_2_U14 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_2_n101), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_2_n105), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_2_n100), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_2_n128) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_2_U13 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_2_n106), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_2_n105) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_2_U12 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_2_n104), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_2_n103) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_2_U11 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_2_n102), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_2_n101) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_2_U10 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_2_n100), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_2_n99) );
  MUX2_X1 SD1_SB_inst_SD1_SB_bit_inst_2_U9 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_2_n97), .B(
        SD1_SB_inst_SD1_SB_bit_inst_2_n98), .S(
        SD1_SB_inst_SD1_SB_bit_inst_2_n99), .Z(
        SD1_SB_inst_SD1_SB_bit_inst_2_n125) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_2_U8 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_2_n118), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_2_n97) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_2_U7 ( .A(CipherErrorVec[4]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_2_n104) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_2_U6 ( .A(CipherErrorVec[2]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_2_n102) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_2_U5 ( .A(CipherErrorVec[5]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_2_n106) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_2_U4 ( .A(CipherErrorVec[1]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_2_n100) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_2_U3 ( .A1(CipherErrorVec[3]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_2_n121), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_2_n98) );
  AOI222_X1 SD1_SB_inst_SD1_SB_bit_inst_3_U45 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_3_n141), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_3_n140), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_3_n141), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_3_n139), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_3_n140), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_3_n138), .ZN(Feedback[63]) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_3_U44 ( .A(StateRegOutput[0]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_3_n137), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_3_n138) );
  AOI211_X1 SD1_SB_inst_SD1_SB_bit_inst_3_U43 ( .C1(
        SD1_SB_inst_SD1_SB_bit_inst_3_n136), .C2(CipherErrorVec[3]), .A(
        SD1_SB_inst_SD1_SB_bit_inst_3_n135), .B(
        SD1_SB_inst_SD1_SB_bit_inst_3_n134), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_3_n137) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_3_U42 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_3_n105), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_3_n103), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_3_n133), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_3_n134) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_3_U41 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_3_n107), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_3_n132), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_3_n131), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_3_n135) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_3_U40 ( .A1(CipherErrorVec[3]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_3_n100), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_3_n131) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_3_U39 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_3_n130), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_3_n136) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_3_U38 ( .A(StateRegOutput[2]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_3_n129), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_3_n139) );
  AOI22_X1 SD1_SB_inst_SD1_SB_bit_inst_3_U37 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_3_n128), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_3_n127), .B1(CipherErrorVec[6]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_3_n126), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_3_n129) );
  OAI211_X1 SD1_SB_inst_SD1_SB_bit_inst_3_U36 ( .C1(
        SD1_SB_inst_SD1_SB_bit_inst_3_n125), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_3_n101), .A(
        SD1_SB_inst_SD1_SB_bit_inst_3_n124), .B(
        SD1_SB_inst_SD1_SB_bit_inst_3_n123), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_3_n126) );
  NAND3_X1 SD1_SB_inst_SD1_SB_bit_inst_3_U35 ( .A1(CipherErrorVec[0]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_3_n108), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_3_n122), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_3_n123) );
  OAI22_X1 SD1_SB_inst_SD1_SB_bit_inst_3_U34 ( .A1(CipherErrorVec[3]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_3_n106), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_3_n100), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_3_n103), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_3_n122) );
  AOI22_X1 SD1_SB_inst_SD1_SB_bit_inst_3_U33 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_3_n102), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_3_n104), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_3_n105), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_3_n108), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_3_n125) );
  OAI21_X1 SD1_SB_inst_SD1_SB_bit_inst_3_U32 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_3_n100), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_3_n121), .A(
        SD1_SB_inst_SD1_SB_bit_inst_3_n120), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_3_n127) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_3_U31 ( .A(CipherErrorVec[0]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_3_n121) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_3_U30 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_3_n124), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_3_n128) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_3_U29 ( .A(StateRegOutput[1]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_3_n119), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_3_n140) );
  AOI22_X1 SD1_SB_inst_SD1_SB_bit_inst_3_U28 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_3_n105), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_3_n118), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_3_n100), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_3_n117), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_3_n119) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_3_U27 ( .A1(CipherErrorVec[3]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_3_n132), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_3_n108), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_3_n117) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_3_U26 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_3_n102), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_3_n105), .A3(CipherErrorVec[0]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_3_n132) );
  OAI22_X1 SD1_SB_inst_SD1_SB_bit_inst_3_U25 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_3_n102), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_3_n133), .B1(CipherErrorVec[6]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_3_n130), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_3_n118) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_3_U24 ( .A1(CipherErrorVec[0]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_3_n116), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_3_n133) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_3_U23 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_3_n115), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_3_n101), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_3_n116) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_3_U22 ( .A1(CipherErrorVec[3]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_3_n107), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_3_n115) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_3_U21 ( .A(StateRegOutput[3]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_3_n114), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_3_n141) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_3_U20 ( .B1(CipherErrorVec[6]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_3_n113), .A(
        SD1_SB_inst_SD1_SB_bit_inst_3_n112), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_3_n114) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_3_U19 ( .B1(CipherErrorVec[0]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_3_n124), .A(
        SD1_SB_inst_SD1_SB_bit_inst_3_n120), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_3_n112) );
  NAND3_X1 SD1_SB_inst_SD1_SB_bit_inst_3_U18 ( .A1(CipherErrorVec[3]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_3_n100), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_3_n107), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_3_n120) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_3_U17 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_3_n102), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_3_n105), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_3_n124) );
  OAI221_X1 SD1_SB_inst_SD1_SB_bit_inst_3_U16 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_3_n105), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_3_n130), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_3_n105), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_3_n111), .A(
        SD1_SB_inst_SD1_SB_bit_inst_3_n110), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_3_n113) );
  OAI21_X1 SD1_SB_inst_SD1_SB_bit_inst_3_U15 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_3_n107), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_3_n109), .A(CipherErrorVec[3]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_3_n110) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_3_U14 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_3_n102), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_3_n100), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_3_n106), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_3_n109) );
  OAI211_X1 SD1_SB_inst_SD1_SB_bit_inst_3_U13 ( .C1(CipherErrorVec[3]), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_3_n107), .A(
        SD1_SB_inst_SD1_SB_bit_inst_3_n100), .B(
        SD1_SB_inst_SD1_SB_bit_inst_3_n103), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_3_n111) );
  NAND3_X1 SD1_SB_inst_SD1_SB_bit_inst_3_U12 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_3_n102), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_3_n107), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_3_n101), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_3_n130) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_3_U11 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_3_n108), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_3_n107) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_3_U10 ( .A(CipherErrorVec[4]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_3_n106) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_3_U9 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_3_n106), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_3_n105) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_3_U8 ( .A(CipherErrorVec[3]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_3_n104) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_3_U7 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_3_n103), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_3_n102) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_3_U6 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_3_n101), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_3_n100) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_3_U5 ( .A(CipherErrorVec[2]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_3_n103) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_3_U4 ( .A(CipherErrorVec[5]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_3_n108) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_3_U3 ( .A(CipherErrorVec[1]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_3_n101) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_4_U47 ( .B1(OutputRegIn[6]), .B2(
        OutputRegIn[7]), .A(SD1_SB_inst_SD1_SB_bit_inst_4_n131), .ZN(
        Feedback[48]) );
  AOI221_X1 SD1_SB_inst_SD1_SB_bit_inst_4_U46 ( .B1(OutputRegIn[6]), .B2(
        OutputRegIn[4]), .C1(OutputRegIn[7]), .C2(OutputRegIn[4]), .A(
        OutputRegIn[5]), .ZN(SD1_SB_inst_SD1_SB_bit_inst_4_n131) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_4_U45 ( .A(StateRegOutput[7]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_4_n127), .ZN(OutputRegIn[7]) );
  AOI211_X1 SD1_SB_inst_SD1_SB_bit_inst_4_U44 ( .C1(CipherErrorVec[13]), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_4_n126), .A(
        SD1_SB_inst_SD1_SB_bit_inst_4_n125), .B(
        SD1_SB_inst_SD1_SB_bit_inst_4_n124), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_4_n127) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_4_U43 ( .A1(CipherErrorVec[7]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_4_n101), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_4_n123), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_4_n124) );
  AOI222_X1 SD1_SB_inst_SD1_SB_bit_inst_4_U42 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_4_n108), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_4_n104), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_4_n108), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_4_n122), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_4_n104), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_4_n121), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_4_n126) );
  OAI221_X1 SD1_SB_inst_SD1_SB_bit_inst_4_U41 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_4_n120), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_4_n100), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_4_n120), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_4_n102), .A(
        SD1_SB_inst_SD1_SB_bit_inst_4_n106), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_4_n121) );
  OAI211_X1 SD1_SB_inst_SD1_SB_bit_inst_4_U40 ( .C1(
        SD1_SB_inst_SD1_SB_bit_inst_4_n105), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_4_n100), .A(
        SD1_SB_inst_SD1_SB_bit_inst_4_n119), .B(
        SD1_SB_inst_SD1_SB_bit_inst_4_n102), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_4_n122) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_4_U39 ( .A(StateRegOutput[6]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_4_n118), .ZN(OutputRegIn[6]) );
  AOI211_X1 SD1_SB_inst_SD1_SB_bit_inst_4_U38 ( .C1(CipherErrorVec[13]), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_4_n117), .A(
        SD1_SB_inst_SD1_SB_bit_inst_4_n125), .B(
        SD1_SB_inst_SD1_SB_bit_inst_4_n116), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_4_n118) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_4_U37 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_4_n128), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_4_n96), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_4_n116) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_4_U36 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_4_n105), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_4_n120), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_4_n128) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_4_U35 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_4_n102), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_4_n123), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_4_n119), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_4_n125) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_4_U34 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_4_n105), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_4_n100), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_4_n119) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_4_U33 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_4_n107), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_4_n103), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_4_n123) );
  OAI22_X1 SD1_SB_inst_SD1_SB_bit_inst_4_U32 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_4_n107), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_4_n115), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_4_n114), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_4_n102), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_4_n117) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_4_U31 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_4_n100), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_4_n104), .A(
        SD1_SB_inst_SD1_SB_bit_inst_4_n105), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_4_n114) );
  AOI22_X1 SD1_SB_inst_SD1_SB_bit_inst_4_U30 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_4_n105), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_4_n100), .B1(CipherErrorVec[7]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_4_n113), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_4_n115) );
  OAI21_X1 SD1_SB_inst_SD1_SB_bit_inst_4_U29 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_4_n103), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_4_n106), .A(
        SD1_SB_inst_SD1_SB_bit_inst_4_n112), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_4_n113) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_4_U28 ( .A(StateRegOutput[4]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_4_n111), .ZN(OutputRegIn[4]) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_4_U27 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_4_n110), .B2(CipherErrorVec[9]), .A(
        SD1_SB_inst_SD1_SB_bit_inst_4_n109), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_4_n111) );
  AOI221_X1 SD1_SB_inst_SD1_SB_bit_inst_4_U26 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_4_n107), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_4_n112), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_4_n108), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_4_n129), .A(
        SD1_SB_inst_SD1_SB_bit_inst_4_n104), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_4_n109) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_4_U25 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_4_n120), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_4_n112) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_4_U24 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_4_n100), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_4_n102), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_4_n120) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_4_U23 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_4_n130), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_4_n105), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_4_n110) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_4_U22 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_4_n108), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_4_n107) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_4_U21 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_4_n106), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_4_n105) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_4_U20 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_4_n104), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_4_n103) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_4_U19 ( .A(CipherErrorVec[9]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_4_n102) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_4_U18 ( .A(CipherErrorVec[8]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_4_n101) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_4_U17 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_4_n101), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_4_n100) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_4_U16 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_4_n99), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_4_n130) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_4_U15 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_4_n97), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_4_n129) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_4_U14 ( .A(CipherErrorVec[7]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_4_n96) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_4_U13 ( .A(CipherErrorVec[12]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_4_n108) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_4_U12 ( .A(CipherErrorVec[11]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_4_n106) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_4_U11 ( .A(CipherErrorVec[10]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_4_n104) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_4_U10 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_4_n100), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_4_n107), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_4_n98) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_4_U9 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_4_n98), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_4_n104), .A(
        SD1_SB_inst_SD1_SB_bit_inst_4_n96), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_4_n99) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_4_U8 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_4_n105), .A2(CipherErrorVec[9]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_4_n95) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_4_U7 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_4_n95), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_4_n96), .A(
        SD1_SB_inst_SD1_SB_bit_inst_4_n101), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_4_n97) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_4_U6 ( .A(StateRegOutput[5]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_4_n94), .ZN(OutputRegIn[5]) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_4_U5 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_4_n107), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_4_n92), .A(
        SD1_SB_inst_SD1_SB_bit_inst_4_n93), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_4_n94) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_4_U4 ( .A1(CipherErrorVec[9]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_4_n130), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_4_n106), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_4_n93) );
  OAI22_X1 SD1_SB_inst_SD1_SB_bit_inst_4_U3 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_4_n103), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_4_n129), .B1(CipherErrorVec[13]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_4_n128), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_4_n92) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_5_U37 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_5_n110), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_5_n109), .A(
        SD1_SB_inst_SD1_SB_bit_inst_5_n108), .ZN(Feedback[49]) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_5_U36 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_5_n107), .B2(StateRegOutput[4]), .A(
        SD1_SB_inst_SD1_SB_bit_inst_5_n106), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_5_n108) );
  OAI22_X1 SD1_SB_inst_SD1_SB_bit_inst_5_U35 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_5_n109), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_5_n110), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_5_n107), .B2(StateRegOutput[4]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_5_n106) );
  AOI22_X1 SD1_SB_inst_SD1_SB_bit_inst_5_U34 ( .A1(CipherErrorVec[7]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_5_n105), .B1(CipherErrorVec[10]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_5_n104), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_5_n107) );
  OAI21_X1 SD1_SB_inst_SD1_SB_bit_inst_5_U33 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_5_n103), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_5_n102), .A(
        SD1_SB_inst_SD1_SB_bit_inst_5_n101), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_5_n104) );
  NAND3_X1 SD1_SB_inst_SD1_SB_bit_inst_5_U32 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_5_n79), .A2(CipherErrorVec[12]), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_5_n78), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_5_n101) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_5_U31 ( .A1(CipherErrorVec[7]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_5_n79), .A3(CipherErrorVec[11]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_5_n103) );
  AOI211_X1 SD1_SB_inst_SD1_SB_bit_inst_5_U30 ( .C1(
        SD1_SB_inst_SD1_SB_bit_inst_5_n100), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_5_n78), .A(CipherErrorVec[11]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_5_n80), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_5_n105) );
  XOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_5_U29 ( .A(StateRegOutput[6]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_5_n99), .Z(
        SD1_SB_inst_SD1_SB_bit_inst_5_n109) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_5_U28 ( .B1(CipherErrorVec[13]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_5_n98), .A(
        SD1_SB_inst_SD1_SB_bit_inst_5_n97), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_5_n99) );
  AOI221_X1 SD1_SB_inst_SD1_SB_bit_inst_5_U27 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_5_n77), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_5_n96), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_5_n78), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_5_n95), .A(
        SD1_SB_inst_SD1_SB_bit_inst_5_n94), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_5_n97) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_5_U26 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_5_n93), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_5_n94) );
  OAI22_X1 SD1_SB_inst_SD1_SB_bit_inst_5_U25 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_5_n92), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_5_n80), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_5_n91), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_5_n82), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_5_n98) );
  AOI211_X1 SD1_SB_inst_SD1_SB_bit_inst_5_U24 ( .C1(CipherErrorVec[7]), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_5_n100), .A(
        SD1_SB_inst_SD1_SB_bit_inst_5_n79), .B(
        SD1_SB_inst_SD1_SB_bit_inst_5_n90), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_5_n91) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_5_U23 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_5_n102), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_5_n90) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_5_U22 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_5_n77), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_5_n83), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_5_n102) );
  AOI22_X1 SD1_SB_inst_SD1_SB_bit_inst_5_U21 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_5_n77), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_5_n81), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_5_n89), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_5_n83), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_5_n92) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_5_U20 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_5_n77), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_5_n95), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_5_n89) );
  XOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_5_U19 ( .A(StateRegOutput[7]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_5_n88), .Z(
        SD1_SB_inst_SD1_SB_bit_inst_5_n110) );
  OAI21_X1 SD1_SB_inst_SD1_SB_bit_inst_5_U18 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_5_n87), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_5_n96), .A(
        SD1_SB_inst_SD1_SB_bit_inst_5_n86), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_5_n88) );
  OAI221_X1 SD1_SB_inst_SD1_SB_bit_inst_5_U17 ( .B1(CipherErrorVec[11]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_5_n85), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_5_n82), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_5_n84), .A(CipherErrorVec[13]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_5_n86) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_5_U16 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_5_n77), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_5_n79), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_5_n81), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_5_n84) );
  OAI33_X1 SD1_SB_inst_SD1_SB_bit_inst_5_U15 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_5_n79), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_5_n100), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_5_n78), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_5_n80), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_5_n83), .B3(
        SD1_SB_inst_SD1_SB_bit_inst_5_n77), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_5_n85) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_5_U14 ( .A1(CipherErrorVec[10]), .A2(
        CipherErrorVec[12]), .ZN(SD1_SB_inst_SD1_SB_bit_inst_5_n100) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_5_U13 ( .A1(CipherErrorVec[10]), .A2(
        CipherErrorVec[12]), .ZN(SD1_SB_inst_SD1_SB_bit_inst_5_n96) );
  AOI221_X1 SD1_SB_inst_SD1_SB_bit_inst_5_U12 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_5_n93), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_5_n77), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_5_n95), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_5_n77), .A(CipherErrorVec[13]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_5_n87) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_5_U11 ( .A(CipherErrorVec[7]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_5_n95) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_5_U10 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_5_n80), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_5_n82), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_5_n93) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_5_U9 ( .A(CipherErrorVec[10]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_5_n81) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_5_U8 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_5_n80), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_5_n79) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_5_U7 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_5_n78), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_5_n77) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_5_U6 ( .A(CipherErrorVec[11]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_5_n82) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_5_U5 ( .A(CipherErrorVec[12]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_5_n83) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_5_U4 ( .A(CipherErrorVec[9]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_5_n80) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_5_U3 ( .A(CipherErrorVec[8]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_5_n78) );
  OAI22_X1 SD1_SB_inst_SD1_SB_bit_inst_6_U45 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_6_n138), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_6_n137), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_6_n136), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_6_n135), .ZN(Feedback[50]) );
  XOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_6_U44 ( .A(StateRegOutput[5]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_6_n134), .Z(
        SD1_SB_inst_SD1_SB_bit_inst_6_n137) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_6_U43 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_6_n103), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_6_n133), .A(
        SD1_SB_inst_SD1_SB_bit_inst_6_n132), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_6_n134) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_6_U42 ( .A1(CipherErrorVec[10]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_6_n131), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_6_n130), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_6_n132) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_6_U41 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_6_n105), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_6_n99), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_6_n130) );
  OAI22_X1 SD1_SB_inst_SD1_SB_bit_inst_6_U40 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_6_n101), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_6_n129), .B1(CipherErrorVec[13]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_6_n128), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_6_n133) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_6_U39 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_6_n135), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_6_n136), .A(
        SD1_SB_inst_SD1_SB_bit_inst_6_n127), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_6_n138) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_6_U38 ( .A(StateRegOutput[6]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_6_n126), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_6_n127) );
  AOI211_X1 SD1_SB_inst_SD1_SB_bit_inst_6_U37 ( .C1(
        SD1_SB_inst_SD1_SB_bit_inst_6_n101), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_6_n125), .A(
        SD1_SB_inst_SD1_SB_bit_inst_6_n124), .B(
        SD1_SB_inst_SD1_SB_bit_inst_6_n123), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_6_n126) );
  AOI211_X1 SD1_SB_inst_SD1_SB_bit_inst_6_U36 ( .C1(
        SD1_SB_inst_SD1_SB_bit_inst_6_n122), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_6_n102), .A(
        SD1_SB_inst_SD1_SB_bit_inst_6_n121), .B(
        SD1_SB_inst_SD1_SB_bit_inst_6_n104), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_6_n123) );
  AOI22_X1 SD1_SB_inst_SD1_SB_bit_inst_6_U35 ( .A1(CipherErrorVec[7]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_6_n120), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_6_n99), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_6_n106), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_6_n122) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_6_U34 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_6_n102), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_6_n104), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_6_n119), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_6_n124) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_6_U33 ( .A(CipherErrorVec[13]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_6_n121) );
  OAI221_X1 SD1_SB_inst_SD1_SB_bit_inst_6_U32 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_6_n103), .B2(CipherErrorVec[13]), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_6_n103), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_6_n106), .A(CipherErrorVec[7]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_6_n118) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_6_U31 ( .A(StateRegOutput[4]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_6_n117), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_6_n136) );
  AOI22_X1 SD1_SB_inst_SD1_SB_bit_inst_6_U30 ( .A1(CipherErrorVec[10]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_6_n116), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_6_n101), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_6_n115), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_6_n117) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_6_U29 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_6_n103), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_6_n129), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_6_n115) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_6_U28 ( .A1(CipherErrorVec[7]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_6_n114), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_6_n129) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_6_U27 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_6_n120), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_6_n100), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_6_n114) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_6_U26 ( .A1(CipherErrorVec[10]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_6_n105), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_6_n120) );
  OAI21_X1 SD1_SB_inst_SD1_SB_bit_inst_6_U25 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_6_n131), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_6_n113), .A(
        SD1_SB_inst_SD1_SB_bit_inst_6_n128), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_6_n116) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_6_U24 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_6_n99), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_6_n106), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_6_n113) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_6_U23 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_6_n101), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_6_n103), .A3(CipherErrorVec[7]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_6_n131) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_6_U22 ( .A(StateRegOutput[7]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_6_n112), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_6_n135) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_6_U21 ( .B1(CipherErrorVec[13]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_6_n111), .A(
        SD1_SB_inst_SD1_SB_bit_inst_6_n110), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_6_n112) );
  AOI221_X1 SD1_SB_inst_SD1_SB_bit_inst_6_U20 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_6_n104), .B2(CipherErrorVec[7]), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_6_n102), .C2(CipherErrorVec[7]), .A(
        SD1_SB_inst_SD1_SB_bit_inst_6_n119), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_6_n110) );
  NAND3_X1 SD1_SB_inst_SD1_SB_bit_inst_6_U19 ( .A1(CipherErrorVec[10]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_6_n105), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_6_n99), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_6_n119) );
  OAI221_X1 SD1_SB_inst_SD1_SB_bit_inst_6_U18 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_6_n103), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_6_n128), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_6_n103), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_6_n109), .A(
        SD1_SB_inst_SD1_SB_bit_inst_6_n108), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_6_n111) );
  OAI21_X1 SD1_SB_inst_SD1_SB_bit_inst_6_U17 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_6_n105), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_6_n107), .A(CipherErrorVec[10]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_6_n108) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_6_U16 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_6_n101), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_6_n99), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_6_n104), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_6_n107) );
  OAI211_X1 SD1_SB_inst_SD1_SB_bit_inst_6_U15 ( .C1(CipherErrorVec[10]), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_6_n105), .A(
        SD1_SB_inst_SD1_SB_bit_inst_6_n99), .B(
        SD1_SB_inst_SD1_SB_bit_inst_6_n102), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_6_n109) );
  NAND3_X1 SD1_SB_inst_SD1_SB_bit_inst_6_U14 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_6_n101), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_6_n105), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_6_n100), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_6_n128) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_6_U13 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_6_n106), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_6_n105) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_6_U12 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_6_n104), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_6_n103) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_6_U11 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_6_n102), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_6_n101) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_6_U10 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_6_n100), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_6_n99) );
  MUX2_X1 SD1_SB_inst_SD1_SB_bit_inst_6_U9 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_6_n97), .B(
        SD1_SB_inst_SD1_SB_bit_inst_6_n98), .S(
        SD1_SB_inst_SD1_SB_bit_inst_6_n99), .Z(
        SD1_SB_inst_SD1_SB_bit_inst_6_n125) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_6_U8 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_6_n118), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_6_n97) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_6_U7 ( .A(CipherErrorVec[11]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_6_n104) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_6_U6 ( .A(CipherErrorVec[9]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_6_n102) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_6_U5 ( .A(CipherErrorVec[12]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_6_n106) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_6_U4 ( .A(CipherErrorVec[8]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_6_n100) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_6_U3 ( .A1(CipherErrorVec[10]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_6_n121), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_6_n98) );
  AOI222_X1 SD1_SB_inst_SD1_SB_bit_inst_7_U45 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_7_n141), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_7_n140), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_7_n141), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_7_n139), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_7_n140), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_7_n138), .ZN(Feedback[51]) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_7_U44 ( .A(StateRegOutput[4]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_7_n137), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_7_n138) );
  AOI211_X1 SD1_SB_inst_SD1_SB_bit_inst_7_U43 ( .C1(
        SD1_SB_inst_SD1_SB_bit_inst_7_n136), .C2(CipherErrorVec[10]), .A(
        SD1_SB_inst_SD1_SB_bit_inst_7_n135), .B(
        SD1_SB_inst_SD1_SB_bit_inst_7_n134), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_7_n137) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_7_U42 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_7_n105), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_7_n103), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_7_n133), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_7_n134) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_7_U41 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_7_n107), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_7_n132), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_7_n131), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_7_n135) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_7_U40 ( .A1(CipherErrorVec[10]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_7_n100), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_7_n131) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_7_U39 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_7_n130), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_7_n136) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_7_U38 ( .A(StateRegOutput[6]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_7_n129), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_7_n139) );
  AOI22_X1 SD1_SB_inst_SD1_SB_bit_inst_7_U37 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_7_n128), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_7_n127), .B1(CipherErrorVec[13]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_7_n126), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_7_n129) );
  OAI211_X1 SD1_SB_inst_SD1_SB_bit_inst_7_U36 ( .C1(
        SD1_SB_inst_SD1_SB_bit_inst_7_n125), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_7_n101), .A(
        SD1_SB_inst_SD1_SB_bit_inst_7_n124), .B(
        SD1_SB_inst_SD1_SB_bit_inst_7_n123), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_7_n126) );
  NAND3_X1 SD1_SB_inst_SD1_SB_bit_inst_7_U35 ( .A1(CipherErrorVec[7]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_7_n108), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_7_n122), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_7_n123) );
  OAI22_X1 SD1_SB_inst_SD1_SB_bit_inst_7_U34 ( .A1(CipherErrorVec[10]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_7_n106), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_7_n100), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_7_n103), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_7_n122) );
  AOI22_X1 SD1_SB_inst_SD1_SB_bit_inst_7_U33 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_7_n102), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_7_n104), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_7_n105), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_7_n108), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_7_n125) );
  OAI21_X1 SD1_SB_inst_SD1_SB_bit_inst_7_U32 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_7_n100), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_7_n121), .A(
        SD1_SB_inst_SD1_SB_bit_inst_7_n120), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_7_n127) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_7_U31 ( .A(CipherErrorVec[7]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_7_n121) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_7_U30 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_7_n124), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_7_n128) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_7_U29 ( .A(StateRegOutput[5]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_7_n119), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_7_n140) );
  AOI22_X1 SD1_SB_inst_SD1_SB_bit_inst_7_U28 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_7_n105), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_7_n118), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_7_n100), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_7_n117), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_7_n119) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_7_U27 ( .A1(CipherErrorVec[10]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_7_n132), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_7_n108), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_7_n117) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_7_U26 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_7_n102), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_7_n105), .A3(CipherErrorVec[7]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_7_n132) );
  OAI22_X1 SD1_SB_inst_SD1_SB_bit_inst_7_U25 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_7_n102), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_7_n133), .B1(CipherErrorVec[13]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_7_n130), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_7_n118) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_7_U24 ( .A1(CipherErrorVec[7]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_7_n116), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_7_n133) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_7_U23 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_7_n115), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_7_n101), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_7_n116) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_7_U22 ( .A1(CipherErrorVec[10]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_7_n107), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_7_n115) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_7_U21 ( .A(StateRegOutput[7]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_7_n114), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_7_n141) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_7_U20 ( .B1(CipherErrorVec[13]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_7_n113), .A(
        SD1_SB_inst_SD1_SB_bit_inst_7_n112), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_7_n114) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_7_U19 ( .B1(CipherErrorVec[7]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_7_n124), .A(
        SD1_SB_inst_SD1_SB_bit_inst_7_n120), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_7_n112) );
  NAND3_X1 SD1_SB_inst_SD1_SB_bit_inst_7_U18 ( .A1(CipherErrorVec[10]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_7_n100), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_7_n107), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_7_n120) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_7_U17 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_7_n102), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_7_n105), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_7_n124) );
  OAI221_X1 SD1_SB_inst_SD1_SB_bit_inst_7_U16 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_7_n105), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_7_n130), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_7_n105), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_7_n111), .A(
        SD1_SB_inst_SD1_SB_bit_inst_7_n110), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_7_n113) );
  OAI21_X1 SD1_SB_inst_SD1_SB_bit_inst_7_U15 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_7_n107), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_7_n109), .A(CipherErrorVec[10]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_7_n110) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_7_U14 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_7_n102), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_7_n100), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_7_n106), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_7_n109) );
  OAI211_X1 SD1_SB_inst_SD1_SB_bit_inst_7_U13 ( .C1(CipherErrorVec[10]), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_7_n107), .A(
        SD1_SB_inst_SD1_SB_bit_inst_7_n100), .B(
        SD1_SB_inst_SD1_SB_bit_inst_7_n103), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_7_n111) );
  NAND3_X1 SD1_SB_inst_SD1_SB_bit_inst_7_U12 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_7_n102), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_7_n107), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_7_n101), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_7_n130) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_7_U11 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_7_n108), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_7_n107) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_7_U10 ( .A(CipherErrorVec[11]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_7_n106) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_7_U9 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_7_n106), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_7_n105) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_7_U8 ( .A(CipherErrorVec[10]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_7_n104) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_7_U7 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_7_n103), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_7_n102) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_7_U6 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_7_n101), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_7_n100) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_7_U5 ( .A(CipherErrorVec[9]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_7_n103) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_7_U4 ( .A(CipherErrorVec[12]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_7_n108) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_7_U3 ( .A(CipherErrorVec[8]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_7_n101) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_8_U47 ( .B1(OutputRegIn[10]), .B2(
        OutputRegIn[11]), .A(SD1_SB_inst_SD1_SB_bit_inst_8_n131), .ZN(
        Feedback[52]) );
  AOI221_X1 SD1_SB_inst_SD1_SB_bit_inst_8_U46 ( .B1(OutputRegIn[10]), .B2(
        OutputRegIn[8]), .C1(OutputRegIn[11]), .C2(OutputRegIn[8]), .A(
        OutputRegIn[9]), .ZN(SD1_SB_inst_SD1_SB_bit_inst_8_n131) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_8_U45 ( .A(StateRegOutput[11]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_8_n127), .ZN(OutputRegIn[11]) );
  AOI211_X1 SD1_SB_inst_SD1_SB_bit_inst_8_U44 ( .C1(CipherErrorVec[20]), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_8_n126), .A(
        SD1_SB_inst_SD1_SB_bit_inst_8_n125), .B(
        SD1_SB_inst_SD1_SB_bit_inst_8_n124), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_8_n127) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_8_U43 ( .A1(CipherErrorVec[14]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_8_n101), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_8_n123), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_8_n124) );
  AOI222_X1 SD1_SB_inst_SD1_SB_bit_inst_8_U42 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_8_n108), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_8_n104), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_8_n108), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_8_n122), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_8_n104), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_8_n121), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_8_n126) );
  OAI221_X1 SD1_SB_inst_SD1_SB_bit_inst_8_U41 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_8_n120), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_8_n100), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_8_n120), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_8_n102), .A(
        SD1_SB_inst_SD1_SB_bit_inst_8_n106), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_8_n121) );
  OAI211_X1 SD1_SB_inst_SD1_SB_bit_inst_8_U40 ( .C1(
        SD1_SB_inst_SD1_SB_bit_inst_8_n105), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_8_n100), .A(
        SD1_SB_inst_SD1_SB_bit_inst_8_n119), .B(
        SD1_SB_inst_SD1_SB_bit_inst_8_n102), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_8_n122) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_8_U39 ( .A(StateRegOutput[10]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_8_n118), .ZN(OutputRegIn[10]) );
  AOI211_X1 SD1_SB_inst_SD1_SB_bit_inst_8_U38 ( .C1(CipherErrorVec[20]), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_8_n117), .A(
        SD1_SB_inst_SD1_SB_bit_inst_8_n125), .B(
        SD1_SB_inst_SD1_SB_bit_inst_8_n116), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_8_n118) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_8_U37 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_8_n128), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_8_n96), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_8_n116) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_8_U36 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_8_n105), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_8_n120), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_8_n128) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_8_U35 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_8_n102), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_8_n123), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_8_n119), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_8_n125) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_8_U34 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_8_n105), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_8_n100), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_8_n119) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_8_U33 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_8_n107), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_8_n103), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_8_n123) );
  OAI22_X1 SD1_SB_inst_SD1_SB_bit_inst_8_U32 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_8_n107), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_8_n115), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_8_n114), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_8_n102), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_8_n117) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_8_U31 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_8_n100), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_8_n104), .A(
        SD1_SB_inst_SD1_SB_bit_inst_8_n105), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_8_n114) );
  AOI22_X1 SD1_SB_inst_SD1_SB_bit_inst_8_U30 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_8_n105), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_8_n100), .B1(CipherErrorVec[14]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_8_n113), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_8_n115) );
  OAI21_X1 SD1_SB_inst_SD1_SB_bit_inst_8_U29 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_8_n103), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_8_n106), .A(
        SD1_SB_inst_SD1_SB_bit_inst_8_n112), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_8_n113) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_8_U28 ( .A(StateRegOutput[8]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_8_n111), .ZN(OutputRegIn[8]) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_8_U27 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_8_n110), .B2(CipherErrorVec[16]), .A(
        SD1_SB_inst_SD1_SB_bit_inst_8_n109), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_8_n111) );
  AOI221_X1 SD1_SB_inst_SD1_SB_bit_inst_8_U26 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_8_n107), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_8_n112), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_8_n108), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_8_n129), .A(
        SD1_SB_inst_SD1_SB_bit_inst_8_n104), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_8_n109) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_8_U25 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_8_n120), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_8_n112) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_8_U24 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_8_n100), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_8_n102), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_8_n120) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_8_U23 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_8_n130), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_8_n105), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_8_n110) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_8_U22 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_8_n108), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_8_n107) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_8_U21 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_8_n106), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_8_n105) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_8_U20 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_8_n104), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_8_n103) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_8_U19 ( .A(CipherErrorVec[16]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_8_n102) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_8_U18 ( .A(CipherErrorVec[15]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_8_n101) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_8_U17 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_8_n101), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_8_n100) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_8_U16 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_8_n99), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_8_n130) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_8_U15 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_8_n97), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_8_n129) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_8_U14 ( .A(CipherErrorVec[14]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_8_n96) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_8_U13 ( .A(CipherErrorVec[19]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_8_n108) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_8_U12 ( .A(CipherErrorVec[18]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_8_n106) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_8_U11 ( .A(CipherErrorVec[17]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_8_n104) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_8_U10 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_8_n100), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_8_n107), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_8_n98) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_8_U9 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_8_n98), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_8_n104), .A(
        SD1_SB_inst_SD1_SB_bit_inst_8_n96), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_8_n99) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_8_U8 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_8_n105), .A2(CipherErrorVec[16]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_8_n95) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_8_U7 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_8_n95), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_8_n96), .A(
        SD1_SB_inst_SD1_SB_bit_inst_8_n101), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_8_n97) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_8_U6 ( .A(StateRegOutput[9]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_8_n94), .ZN(OutputRegIn[9]) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_8_U5 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_8_n107), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_8_n92), .A(
        SD1_SB_inst_SD1_SB_bit_inst_8_n93), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_8_n94) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_8_U4 ( .A1(CipherErrorVec[16]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_8_n130), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_8_n106), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_8_n93) );
  OAI22_X1 SD1_SB_inst_SD1_SB_bit_inst_8_U3 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_8_n103), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_8_n129), .B1(CipherErrorVec[20]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_8_n128), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_8_n92) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_9_U37 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_9_n110), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_9_n109), .A(
        SD1_SB_inst_SD1_SB_bit_inst_9_n108), .ZN(Feedback[53]) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_9_U36 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_9_n107), .B2(StateRegOutput[8]), .A(
        SD1_SB_inst_SD1_SB_bit_inst_9_n106), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_9_n108) );
  OAI22_X1 SD1_SB_inst_SD1_SB_bit_inst_9_U35 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_9_n109), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_9_n110), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_9_n107), .B2(StateRegOutput[8]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_9_n106) );
  AOI22_X1 SD1_SB_inst_SD1_SB_bit_inst_9_U34 ( .A1(CipherErrorVec[14]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_9_n105), .B1(CipherErrorVec[17]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_9_n104), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_9_n107) );
  OAI21_X1 SD1_SB_inst_SD1_SB_bit_inst_9_U33 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_9_n103), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_9_n102), .A(
        SD1_SB_inst_SD1_SB_bit_inst_9_n101), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_9_n104) );
  NAND3_X1 SD1_SB_inst_SD1_SB_bit_inst_9_U32 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_9_n79), .A2(CipherErrorVec[19]), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_9_n78), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_9_n101) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_9_U31 ( .A1(CipherErrorVec[14]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_9_n79), .A3(CipherErrorVec[18]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_9_n103) );
  AOI211_X1 SD1_SB_inst_SD1_SB_bit_inst_9_U30 ( .C1(
        SD1_SB_inst_SD1_SB_bit_inst_9_n100), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_9_n78), .A(CipherErrorVec[18]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_9_n80), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_9_n105) );
  XOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_9_U29 ( .A(StateRegOutput[10]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_9_n99), .Z(
        SD1_SB_inst_SD1_SB_bit_inst_9_n109) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_9_U28 ( .B1(CipherErrorVec[20]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_9_n98), .A(
        SD1_SB_inst_SD1_SB_bit_inst_9_n97), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_9_n99) );
  AOI221_X1 SD1_SB_inst_SD1_SB_bit_inst_9_U27 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_9_n77), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_9_n96), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_9_n78), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_9_n95), .A(
        SD1_SB_inst_SD1_SB_bit_inst_9_n94), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_9_n97) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_9_U26 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_9_n93), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_9_n94) );
  OAI22_X1 SD1_SB_inst_SD1_SB_bit_inst_9_U25 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_9_n92), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_9_n80), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_9_n91), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_9_n82), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_9_n98) );
  AOI211_X1 SD1_SB_inst_SD1_SB_bit_inst_9_U24 ( .C1(CipherErrorVec[14]), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_9_n100), .A(
        SD1_SB_inst_SD1_SB_bit_inst_9_n79), .B(
        SD1_SB_inst_SD1_SB_bit_inst_9_n90), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_9_n91) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_9_U23 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_9_n102), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_9_n90) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_9_U22 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_9_n77), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_9_n83), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_9_n102) );
  AOI22_X1 SD1_SB_inst_SD1_SB_bit_inst_9_U21 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_9_n77), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_9_n81), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_9_n89), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_9_n83), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_9_n92) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_9_U20 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_9_n77), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_9_n95), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_9_n89) );
  XOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_9_U19 ( .A(StateRegOutput[11]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_9_n88), .Z(
        SD1_SB_inst_SD1_SB_bit_inst_9_n110) );
  OAI21_X1 SD1_SB_inst_SD1_SB_bit_inst_9_U18 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_9_n87), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_9_n96), .A(
        SD1_SB_inst_SD1_SB_bit_inst_9_n86), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_9_n88) );
  OAI221_X1 SD1_SB_inst_SD1_SB_bit_inst_9_U17 ( .B1(CipherErrorVec[18]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_9_n85), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_9_n82), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_9_n84), .A(CipherErrorVec[20]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_9_n86) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_9_U16 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_9_n77), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_9_n79), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_9_n81), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_9_n84) );
  OAI33_X1 SD1_SB_inst_SD1_SB_bit_inst_9_U15 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_9_n79), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_9_n100), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_9_n78), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_9_n80), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_9_n83), .B3(
        SD1_SB_inst_SD1_SB_bit_inst_9_n77), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_9_n85) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_9_U14 ( .A1(CipherErrorVec[17]), .A2(
        CipherErrorVec[19]), .ZN(SD1_SB_inst_SD1_SB_bit_inst_9_n100) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_9_U13 ( .A1(CipherErrorVec[17]), .A2(
        CipherErrorVec[19]), .ZN(SD1_SB_inst_SD1_SB_bit_inst_9_n96) );
  AOI221_X1 SD1_SB_inst_SD1_SB_bit_inst_9_U12 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_9_n93), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_9_n77), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_9_n95), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_9_n77), .A(CipherErrorVec[20]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_9_n87) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_9_U11 ( .A(CipherErrorVec[14]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_9_n95) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_9_U10 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_9_n80), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_9_n82), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_9_n93) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_9_U9 ( .A(CipherErrorVec[17]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_9_n81) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_9_U8 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_9_n80), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_9_n79) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_9_U7 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_9_n78), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_9_n77) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_9_U6 ( .A(CipherErrorVec[18]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_9_n82) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_9_U5 ( .A(CipherErrorVec[19]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_9_n83) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_9_U4 ( .A(CipherErrorVec[16]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_9_n80) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_9_U3 ( .A(CipherErrorVec[15]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_9_n78) );
  OAI22_X1 SD1_SB_inst_SD1_SB_bit_inst_10_U45 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_10_n138), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_10_n137), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_10_n136), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_10_n135), .ZN(Feedback[54]) );
  XOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_10_U44 ( .A(StateRegOutput[9]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_10_n134), .Z(
        SD1_SB_inst_SD1_SB_bit_inst_10_n137) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_10_U43 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_10_n103), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_10_n133), .A(
        SD1_SB_inst_SD1_SB_bit_inst_10_n132), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_10_n134) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_10_U42 ( .A1(CipherErrorVec[17]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_10_n131), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_10_n130), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_10_n132) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_10_U41 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_10_n105), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_10_n99), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_10_n130) );
  OAI22_X1 SD1_SB_inst_SD1_SB_bit_inst_10_U40 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_10_n101), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_10_n129), .B1(CipherErrorVec[20]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_10_n128), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_10_n133) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_10_U39 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_10_n135), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_10_n136), .A(
        SD1_SB_inst_SD1_SB_bit_inst_10_n127), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_10_n138) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_10_U38 ( .A(StateRegOutput[10]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_10_n126), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_10_n127) );
  AOI211_X1 SD1_SB_inst_SD1_SB_bit_inst_10_U37 ( .C1(
        SD1_SB_inst_SD1_SB_bit_inst_10_n101), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_10_n125), .A(
        SD1_SB_inst_SD1_SB_bit_inst_10_n124), .B(
        SD1_SB_inst_SD1_SB_bit_inst_10_n123), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_10_n126) );
  AOI211_X1 SD1_SB_inst_SD1_SB_bit_inst_10_U36 ( .C1(
        SD1_SB_inst_SD1_SB_bit_inst_10_n122), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_10_n102), .A(
        SD1_SB_inst_SD1_SB_bit_inst_10_n121), .B(
        SD1_SB_inst_SD1_SB_bit_inst_10_n104), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_10_n123) );
  AOI22_X1 SD1_SB_inst_SD1_SB_bit_inst_10_U35 ( .A1(CipherErrorVec[14]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_10_n120), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_10_n99), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_10_n106), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_10_n122) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_10_U34 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_10_n102), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_10_n104), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_10_n119), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_10_n124) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_10_U33 ( .A(CipherErrorVec[20]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_10_n121) );
  OAI221_X1 SD1_SB_inst_SD1_SB_bit_inst_10_U32 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_10_n103), .B2(CipherErrorVec[20]), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_10_n103), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_10_n106), .A(CipherErrorVec[14]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_10_n118) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_10_U31 ( .A(StateRegOutput[8]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_10_n117), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_10_n136) );
  AOI22_X1 SD1_SB_inst_SD1_SB_bit_inst_10_U30 ( .A1(CipherErrorVec[17]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_10_n116), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_10_n101), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_10_n115), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_10_n117) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_10_U29 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_10_n103), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_10_n129), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_10_n115) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_10_U28 ( .A1(CipherErrorVec[14]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_10_n114), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_10_n129) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_10_U27 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_10_n120), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_10_n100), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_10_n114) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_10_U26 ( .A1(CipherErrorVec[17]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_10_n105), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_10_n120) );
  OAI21_X1 SD1_SB_inst_SD1_SB_bit_inst_10_U25 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_10_n131), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_10_n113), .A(
        SD1_SB_inst_SD1_SB_bit_inst_10_n128), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_10_n116) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_10_U24 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_10_n99), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_10_n106), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_10_n113) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_10_U23 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_10_n101), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_10_n103), .A3(CipherErrorVec[14]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_10_n131) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_10_U22 ( .A(StateRegOutput[11]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_10_n112), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_10_n135) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_10_U21 ( .B1(CipherErrorVec[20]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_10_n111), .A(
        SD1_SB_inst_SD1_SB_bit_inst_10_n110), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_10_n112) );
  AOI221_X1 SD1_SB_inst_SD1_SB_bit_inst_10_U20 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_10_n104), .B2(CipherErrorVec[14]), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_10_n102), .C2(CipherErrorVec[14]), .A(
        SD1_SB_inst_SD1_SB_bit_inst_10_n119), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_10_n110) );
  NAND3_X1 SD1_SB_inst_SD1_SB_bit_inst_10_U19 ( .A1(CipherErrorVec[17]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_10_n105), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_10_n99), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_10_n119) );
  OAI221_X1 SD1_SB_inst_SD1_SB_bit_inst_10_U18 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_10_n103), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_10_n128), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_10_n103), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_10_n109), .A(
        SD1_SB_inst_SD1_SB_bit_inst_10_n108), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_10_n111) );
  OAI21_X1 SD1_SB_inst_SD1_SB_bit_inst_10_U17 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_10_n105), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_10_n107), .A(CipherErrorVec[17]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_10_n108) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_10_U16 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_10_n101), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_10_n99), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_10_n104), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_10_n107) );
  OAI211_X1 SD1_SB_inst_SD1_SB_bit_inst_10_U15 ( .C1(CipherErrorVec[17]), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_10_n105), .A(
        SD1_SB_inst_SD1_SB_bit_inst_10_n99), .B(
        SD1_SB_inst_SD1_SB_bit_inst_10_n102), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_10_n109) );
  NAND3_X1 SD1_SB_inst_SD1_SB_bit_inst_10_U14 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_10_n101), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_10_n105), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_10_n100), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_10_n128) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_10_U13 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_10_n106), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_10_n105) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_10_U12 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_10_n104), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_10_n103) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_10_U11 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_10_n102), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_10_n101) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_10_U10 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_10_n100), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_10_n99) );
  MUX2_X1 SD1_SB_inst_SD1_SB_bit_inst_10_U9 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_10_n97), .B(
        SD1_SB_inst_SD1_SB_bit_inst_10_n98), .S(
        SD1_SB_inst_SD1_SB_bit_inst_10_n99), .Z(
        SD1_SB_inst_SD1_SB_bit_inst_10_n125) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_10_U8 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_10_n118), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_10_n97) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_10_U7 ( .A(CipherErrorVec[18]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_10_n104) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_10_U6 ( .A(CipherErrorVec[16]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_10_n102) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_10_U5 ( .A(CipherErrorVec[19]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_10_n106) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_10_U4 ( .A(CipherErrorVec[15]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_10_n100) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_10_U3 ( .A1(CipherErrorVec[17]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_10_n121), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_10_n98) );
  AOI222_X1 SD1_SB_inst_SD1_SB_bit_inst_11_U45 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_11_n141), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_11_n140), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_11_n141), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_11_n139), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_11_n140), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_11_n138), .ZN(Feedback[55]) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_11_U44 ( .A(StateRegOutput[8]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_11_n137), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_11_n138) );
  AOI211_X1 SD1_SB_inst_SD1_SB_bit_inst_11_U43 ( .C1(
        SD1_SB_inst_SD1_SB_bit_inst_11_n136), .C2(CipherErrorVec[17]), .A(
        SD1_SB_inst_SD1_SB_bit_inst_11_n135), .B(
        SD1_SB_inst_SD1_SB_bit_inst_11_n134), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_11_n137) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_11_U42 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_11_n105), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_11_n103), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_11_n133), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_11_n134) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_11_U41 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_11_n107), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_11_n132), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_11_n131), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_11_n135) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_11_U40 ( .A1(CipherErrorVec[17]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_11_n100), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_11_n131) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_11_U39 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_11_n130), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_11_n136) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_11_U38 ( .A(StateRegOutput[10]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_11_n129), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_11_n139) );
  AOI22_X1 SD1_SB_inst_SD1_SB_bit_inst_11_U37 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_11_n128), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_11_n127), .B1(CipherErrorVec[20]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_11_n126), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_11_n129) );
  OAI211_X1 SD1_SB_inst_SD1_SB_bit_inst_11_U36 ( .C1(
        SD1_SB_inst_SD1_SB_bit_inst_11_n125), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_11_n101), .A(
        SD1_SB_inst_SD1_SB_bit_inst_11_n124), .B(
        SD1_SB_inst_SD1_SB_bit_inst_11_n123), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_11_n126) );
  NAND3_X1 SD1_SB_inst_SD1_SB_bit_inst_11_U35 ( .A1(CipherErrorVec[14]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_11_n108), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_11_n122), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_11_n123) );
  OAI22_X1 SD1_SB_inst_SD1_SB_bit_inst_11_U34 ( .A1(CipherErrorVec[17]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_11_n106), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_11_n100), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_11_n103), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_11_n122) );
  AOI22_X1 SD1_SB_inst_SD1_SB_bit_inst_11_U33 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_11_n102), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_11_n104), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_11_n105), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_11_n108), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_11_n125) );
  OAI21_X1 SD1_SB_inst_SD1_SB_bit_inst_11_U32 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_11_n100), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_11_n121), .A(
        SD1_SB_inst_SD1_SB_bit_inst_11_n120), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_11_n127) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_11_U31 ( .A(CipherErrorVec[14]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_11_n121) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_11_U30 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_11_n124), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_11_n128) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_11_U29 ( .A(StateRegOutput[9]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_11_n119), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_11_n140) );
  AOI22_X1 SD1_SB_inst_SD1_SB_bit_inst_11_U28 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_11_n105), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_11_n118), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_11_n100), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_11_n117), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_11_n119) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_11_U27 ( .A1(CipherErrorVec[17]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_11_n132), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_11_n108), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_11_n117) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_11_U26 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_11_n102), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_11_n105), .A3(CipherErrorVec[14]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_11_n132) );
  OAI22_X1 SD1_SB_inst_SD1_SB_bit_inst_11_U25 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_11_n102), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_11_n133), .B1(CipherErrorVec[20]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_11_n130), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_11_n118) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_11_U24 ( .A1(CipherErrorVec[14]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_11_n116), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_11_n133) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_11_U23 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_11_n115), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_11_n101), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_11_n116) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_11_U22 ( .A1(CipherErrorVec[17]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_11_n107), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_11_n115) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_11_U21 ( .A(StateRegOutput[11]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_11_n114), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_11_n141) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_11_U20 ( .B1(CipherErrorVec[20]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_11_n113), .A(
        SD1_SB_inst_SD1_SB_bit_inst_11_n112), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_11_n114) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_11_U19 ( .B1(CipherErrorVec[14]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_11_n124), .A(
        SD1_SB_inst_SD1_SB_bit_inst_11_n120), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_11_n112) );
  NAND3_X1 SD1_SB_inst_SD1_SB_bit_inst_11_U18 ( .A1(CipherErrorVec[17]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_11_n100), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_11_n107), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_11_n120) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_11_U17 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_11_n102), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_11_n105), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_11_n124) );
  OAI221_X1 SD1_SB_inst_SD1_SB_bit_inst_11_U16 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_11_n105), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_11_n130), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_11_n105), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_11_n111), .A(
        SD1_SB_inst_SD1_SB_bit_inst_11_n110), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_11_n113) );
  OAI21_X1 SD1_SB_inst_SD1_SB_bit_inst_11_U15 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_11_n107), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_11_n109), .A(CipherErrorVec[17]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_11_n110) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_11_U14 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_11_n102), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_11_n100), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_11_n106), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_11_n109) );
  OAI211_X1 SD1_SB_inst_SD1_SB_bit_inst_11_U13 ( .C1(CipherErrorVec[17]), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_11_n107), .A(
        SD1_SB_inst_SD1_SB_bit_inst_11_n100), .B(
        SD1_SB_inst_SD1_SB_bit_inst_11_n103), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_11_n111) );
  NAND3_X1 SD1_SB_inst_SD1_SB_bit_inst_11_U12 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_11_n102), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_11_n107), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_11_n101), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_11_n130) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_11_U11 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_11_n108), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_11_n107) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_11_U10 ( .A(CipherErrorVec[18]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_11_n106) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_11_U9 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_11_n106), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_11_n105) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_11_U8 ( .A(CipherErrorVec[17]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_11_n104) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_11_U7 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_11_n103), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_11_n102) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_11_U6 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_11_n101), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_11_n100) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_11_U5 ( .A(CipherErrorVec[16]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_11_n103) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_11_U4 ( .A(CipherErrorVec[19]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_11_n108) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_11_U3 ( .A(CipherErrorVec[15]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_11_n101) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_12_U47 ( .B1(OutputRegIn[14]), .B2(
        OutputRegIn[15]), .A(SD1_SB_inst_SD1_SB_bit_inst_12_n131), .ZN(
        Feedback[56]) );
  AOI221_X1 SD1_SB_inst_SD1_SB_bit_inst_12_U46 ( .B1(OutputRegIn[14]), .B2(
        OutputRegIn[12]), .C1(OutputRegIn[15]), .C2(OutputRegIn[12]), .A(
        OutputRegIn[13]), .ZN(SD1_SB_inst_SD1_SB_bit_inst_12_n131) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_12_U45 ( .A(StateRegOutput[15]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_12_n127), .ZN(OutputRegIn[15]) );
  AOI211_X1 SD1_SB_inst_SD1_SB_bit_inst_12_U44 ( .C1(CipherErrorVec[27]), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_12_n126), .A(
        SD1_SB_inst_SD1_SB_bit_inst_12_n125), .B(
        SD1_SB_inst_SD1_SB_bit_inst_12_n124), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_12_n127) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_12_U43 ( .A1(CipherErrorVec[21]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_12_n101), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_12_n123), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_12_n124) );
  AOI222_X1 SD1_SB_inst_SD1_SB_bit_inst_12_U42 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_12_n108), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_12_n104), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_12_n108), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_12_n122), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_12_n104), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_12_n121), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_12_n126) );
  OAI221_X1 SD1_SB_inst_SD1_SB_bit_inst_12_U41 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_12_n120), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_12_n100), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_12_n120), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_12_n102), .A(
        SD1_SB_inst_SD1_SB_bit_inst_12_n106), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_12_n121) );
  OAI211_X1 SD1_SB_inst_SD1_SB_bit_inst_12_U40 ( .C1(
        SD1_SB_inst_SD1_SB_bit_inst_12_n105), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_12_n100), .A(
        SD1_SB_inst_SD1_SB_bit_inst_12_n119), .B(
        SD1_SB_inst_SD1_SB_bit_inst_12_n102), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_12_n122) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_12_U39 ( .A(StateRegOutput[14]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_12_n118), .ZN(OutputRegIn[14]) );
  AOI211_X1 SD1_SB_inst_SD1_SB_bit_inst_12_U38 ( .C1(CipherErrorVec[27]), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_12_n117), .A(
        SD1_SB_inst_SD1_SB_bit_inst_12_n125), .B(
        SD1_SB_inst_SD1_SB_bit_inst_12_n116), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_12_n118) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_12_U37 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_12_n128), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_12_n96), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_12_n116) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_12_U36 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_12_n105), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_12_n120), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_12_n128) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_12_U35 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_12_n102), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_12_n123), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_12_n119), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_12_n125) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_12_U34 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_12_n105), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_12_n100), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_12_n119) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_12_U33 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_12_n107), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_12_n103), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_12_n123) );
  OAI22_X1 SD1_SB_inst_SD1_SB_bit_inst_12_U32 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_12_n107), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_12_n115), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_12_n114), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_12_n102), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_12_n117) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_12_U31 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_12_n100), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_12_n104), .A(
        SD1_SB_inst_SD1_SB_bit_inst_12_n105), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_12_n114) );
  AOI22_X1 SD1_SB_inst_SD1_SB_bit_inst_12_U30 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_12_n105), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_12_n100), .B1(CipherErrorVec[21]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_12_n113), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_12_n115) );
  OAI21_X1 SD1_SB_inst_SD1_SB_bit_inst_12_U29 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_12_n103), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_12_n106), .A(
        SD1_SB_inst_SD1_SB_bit_inst_12_n112), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_12_n113) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_12_U28 ( .A(StateRegOutput[12]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_12_n111), .ZN(OutputRegIn[12]) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_12_U27 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_12_n110), .B2(CipherErrorVec[23]), .A(
        SD1_SB_inst_SD1_SB_bit_inst_12_n109), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_12_n111) );
  AOI221_X1 SD1_SB_inst_SD1_SB_bit_inst_12_U26 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_12_n107), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_12_n112), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_12_n108), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_12_n129), .A(
        SD1_SB_inst_SD1_SB_bit_inst_12_n104), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_12_n109) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_12_U25 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_12_n120), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_12_n112) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_12_U24 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_12_n100), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_12_n102), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_12_n120) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_12_U23 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_12_n130), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_12_n105), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_12_n110) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_12_U22 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_12_n108), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_12_n107) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_12_U21 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_12_n106), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_12_n105) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_12_U20 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_12_n104), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_12_n103) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_12_U19 ( .A(CipherErrorVec[23]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_12_n102) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_12_U18 ( .A(CipherErrorVec[22]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_12_n101) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_12_U17 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_12_n101), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_12_n100) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_12_U16 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_12_n99), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_12_n130) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_12_U15 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_12_n97), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_12_n129) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_12_U14 ( .A(CipherErrorVec[21]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_12_n96) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_12_U13 ( .A(CipherErrorVec[26]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_12_n108) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_12_U12 ( .A(CipherErrorVec[25]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_12_n106) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_12_U11 ( .A(CipherErrorVec[24]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_12_n104) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_12_U10 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_12_n100), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_12_n107), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_12_n98) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_12_U9 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_12_n98), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_12_n104), .A(
        SD1_SB_inst_SD1_SB_bit_inst_12_n96), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_12_n99) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_12_U8 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_12_n105), .A2(CipherErrorVec[23]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_12_n95) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_12_U7 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_12_n95), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_12_n96), .A(
        SD1_SB_inst_SD1_SB_bit_inst_12_n101), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_12_n97) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_12_U6 ( .A(StateRegOutput[13]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_12_n94), .ZN(OutputRegIn[13]) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_12_U5 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_12_n107), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_12_n92), .A(
        SD1_SB_inst_SD1_SB_bit_inst_12_n93), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_12_n94) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_12_U4 ( .A1(CipherErrorVec[23]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_12_n130), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_12_n106), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_12_n93) );
  OAI22_X1 SD1_SB_inst_SD1_SB_bit_inst_12_U3 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_12_n103), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_12_n129), .B1(CipherErrorVec[27]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_12_n128), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_12_n92) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_13_U37 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_13_n110), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_13_n109), .A(
        SD1_SB_inst_SD1_SB_bit_inst_13_n108), .ZN(Feedback[57]) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_13_U36 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_13_n107), .B2(StateRegOutput[12]), .A(
        SD1_SB_inst_SD1_SB_bit_inst_13_n106), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_13_n108) );
  OAI22_X1 SD1_SB_inst_SD1_SB_bit_inst_13_U35 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_13_n109), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_13_n110), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_13_n107), .B2(StateRegOutput[12]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_13_n106) );
  AOI22_X1 SD1_SB_inst_SD1_SB_bit_inst_13_U34 ( .A1(CipherErrorVec[21]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_13_n105), .B1(CipherErrorVec[24]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_13_n104), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_13_n107) );
  OAI21_X1 SD1_SB_inst_SD1_SB_bit_inst_13_U33 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_13_n103), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_13_n102), .A(
        SD1_SB_inst_SD1_SB_bit_inst_13_n101), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_13_n104) );
  NAND3_X1 SD1_SB_inst_SD1_SB_bit_inst_13_U32 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_13_n79), .A2(CipherErrorVec[26]), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_13_n78), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_13_n101) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_13_U31 ( .A1(CipherErrorVec[21]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_13_n79), .A3(CipherErrorVec[25]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_13_n103) );
  AOI211_X1 SD1_SB_inst_SD1_SB_bit_inst_13_U30 ( .C1(
        SD1_SB_inst_SD1_SB_bit_inst_13_n100), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_13_n78), .A(CipherErrorVec[25]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_13_n80), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_13_n105) );
  XOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_13_U29 ( .A(StateRegOutput[14]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_13_n99), .Z(
        SD1_SB_inst_SD1_SB_bit_inst_13_n109) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_13_U28 ( .B1(CipherErrorVec[27]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_13_n98), .A(
        SD1_SB_inst_SD1_SB_bit_inst_13_n97), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_13_n99) );
  AOI221_X1 SD1_SB_inst_SD1_SB_bit_inst_13_U27 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_13_n77), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_13_n96), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_13_n78), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_13_n95), .A(
        SD1_SB_inst_SD1_SB_bit_inst_13_n94), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_13_n97) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_13_U26 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_13_n93), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_13_n94) );
  OAI22_X1 SD1_SB_inst_SD1_SB_bit_inst_13_U25 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_13_n92), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_13_n80), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_13_n91), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_13_n82), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_13_n98) );
  AOI211_X1 SD1_SB_inst_SD1_SB_bit_inst_13_U24 ( .C1(CipherErrorVec[21]), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_13_n100), .A(
        SD1_SB_inst_SD1_SB_bit_inst_13_n79), .B(
        SD1_SB_inst_SD1_SB_bit_inst_13_n90), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_13_n91) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_13_U23 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_13_n102), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_13_n90) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_13_U22 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_13_n77), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_13_n83), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_13_n102) );
  AOI22_X1 SD1_SB_inst_SD1_SB_bit_inst_13_U21 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_13_n77), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_13_n81), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_13_n89), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_13_n83), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_13_n92) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_13_U20 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_13_n77), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_13_n95), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_13_n89) );
  XOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_13_U19 ( .A(StateRegOutput[15]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_13_n88), .Z(
        SD1_SB_inst_SD1_SB_bit_inst_13_n110) );
  OAI21_X1 SD1_SB_inst_SD1_SB_bit_inst_13_U18 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_13_n87), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_13_n96), .A(
        SD1_SB_inst_SD1_SB_bit_inst_13_n86), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_13_n88) );
  OAI221_X1 SD1_SB_inst_SD1_SB_bit_inst_13_U17 ( .B1(CipherErrorVec[25]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_13_n85), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_13_n82), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_13_n84), .A(CipherErrorVec[27]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_13_n86) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_13_U16 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_13_n77), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_13_n79), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_13_n81), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_13_n84) );
  OAI33_X1 SD1_SB_inst_SD1_SB_bit_inst_13_U15 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_13_n79), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_13_n100), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_13_n78), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_13_n80), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_13_n83), .B3(
        SD1_SB_inst_SD1_SB_bit_inst_13_n77), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_13_n85) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_13_U14 ( .A1(CipherErrorVec[24]), .A2(
        CipherErrorVec[26]), .ZN(SD1_SB_inst_SD1_SB_bit_inst_13_n100) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_13_U13 ( .A1(CipherErrorVec[24]), .A2(
        CipherErrorVec[26]), .ZN(SD1_SB_inst_SD1_SB_bit_inst_13_n96) );
  AOI221_X1 SD1_SB_inst_SD1_SB_bit_inst_13_U12 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_13_n93), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_13_n77), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_13_n95), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_13_n77), .A(CipherErrorVec[27]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_13_n87) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_13_U11 ( .A(CipherErrorVec[21]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_13_n95) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_13_U10 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_13_n80), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_13_n82), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_13_n93) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_13_U9 ( .A(CipherErrorVec[24]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_13_n81) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_13_U8 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_13_n80), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_13_n79) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_13_U7 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_13_n78), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_13_n77) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_13_U6 ( .A(CipherErrorVec[25]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_13_n82) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_13_U5 ( .A(CipherErrorVec[26]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_13_n83) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_13_U4 ( .A(CipherErrorVec[23]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_13_n80) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_13_U3 ( .A(CipherErrorVec[22]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_13_n78) );
  OAI22_X1 SD1_SB_inst_SD1_SB_bit_inst_14_U45 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_14_n138), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_14_n137), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_14_n136), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_14_n135), .ZN(Feedback[58]) );
  XOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_14_U44 ( .A(StateRegOutput[13]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_14_n134), .Z(
        SD1_SB_inst_SD1_SB_bit_inst_14_n137) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_14_U43 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_14_n103), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_14_n133), .A(
        SD1_SB_inst_SD1_SB_bit_inst_14_n132), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_14_n134) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_14_U42 ( .A1(CipherErrorVec[24]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_14_n131), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_14_n130), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_14_n132) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_14_U41 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_14_n105), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_14_n99), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_14_n130) );
  OAI22_X1 SD1_SB_inst_SD1_SB_bit_inst_14_U40 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_14_n101), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_14_n129), .B1(CipherErrorVec[27]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_14_n128), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_14_n133) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_14_U39 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_14_n135), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_14_n136), .A(
        SD1_SB_inst_SD1_SB_bit_inst_14_n127), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_14_n138) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_14_U38 ( .A(StateRegOutput[14]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_14_n126), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_14_n127) );
  AOI211_X1 SD1_SB_inst_SD1_SB_bit_inst_14_U37 ( .C1(
        SD1_SB_inst_SD1_SB_bit_inst_14_n101), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_14_n125), .A(
        SD1_SB_inst_SD1_SB_bit_inst_14_n124), .B(
        SD1_SB_inst_SD1_SB_bit_inst_14_n123), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_14_n126) );
  AOI211_X1 SD1_SB_inst_SD1_SB_bit_inst_14_U36 ( .C1(
        SD1_SB_inst_SD1_SB_bit_inst_14_n122), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_14_n102), .A(
        SD1_SB_inst_SD1_SB_bit_inst_14_n121), .B(
        SD1_SB_inst_SD1_SB_bit_inst_14_n104), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_14_n123) );
  AOI22_X1 SD1_SB_inst_SD1_SB_bit_inst_14_U35 ( .A1(CipherErrorVec[21]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_14_n120), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_14_n99), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_14_n106), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_14_n122) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_14_U34 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_14_n102), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_14_n104), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_14_n119), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_14_n124) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_14_U33 ( .A(CipherErrorVec[27]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_14_n121) );
  OAI221_X1 SD1_SB_inst_SD1_SB_bit_inst_14_U32 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_14_n103), .B2(CipherErrorVec[27]), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_14_n103), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_14_n106), .A(CipherErrorVec[21]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_14_n118) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_14_U31 ( .A(StateRegOutput[12]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_14_n117), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_14_n136) );
  AOI22_X1 SD1_SB_inst_SD1_SB_bit_inst_14_U30 ( .A1(CipherErrorVec[24]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_14_n116), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_14_n101), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_14_n115), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_14_n117) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_14_U29 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_14_n103), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_14_n129), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_14_n115) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_14_U28 ( .A1(CipherErrorVec[21]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_14_n114), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_14_n129) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_14_U27 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_14_n120), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_14_n100), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_14_n114) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_14_U26 ( .A1(CipherErrorVec[24]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_14_n105), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_14_n120) );
  OAI21_X1 SD1_SB_inst_SD1_SB_bit_inst_14_U25 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_14_n131), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_14_n113), .A(
        SD1_SB_inst_SD1_SB_bit_inst_14_n128), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_14_n116) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_14_U24 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_14_n99), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_14_n106), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_14_n113) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_14_U23 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_14_n101), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_14_n103), .A3(CipherErrorVec[21]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_14_n131) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_14_U22 ( .A(StateRegOutput[15]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_14_n112), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_14_n135) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_14_U21 ( .B1(CipherErrorVec[27]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_14_n111), .A(
        SD1_SB_inst_SD1_SB_bit_inst_14_n110), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_14_n112) );
  AOI221_X1 SD1_SB_inst_SD1_SB_bit_inst_14_U20 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_14_n104), .B2(CipherErrorVec[21]), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_14_n102), .C2(CipherErrorVec[21]), .A(
        SD1_SB_inst_SD1_SB_bit_inst_14_n119), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_14_n110) );
  NAND3_X1 SD1_SB_inst_SD1_SB_bit_inst_14_U19 ( .A1(CipherErrorVec[24]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_14_n105), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_14_n99), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_14_n119) );
  OAI221_X1 SD1_SB_inst_SD1_SB_bit_inst_14_U18 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_14_n103), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_14_n128), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_14_n103), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_14_n109), .A(
        SD1_SB_inst_SD1_SB_bit_inst_14_n108), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_14_n111) );
  OAI21_X1 SD1_SB_inst_SD1_SB_bit_inst_14_U17 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_14_n105), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_14_n107), .A(CipherErrorVec[24]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_14_n108) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_14_U16 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_14_n101), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_14_n99), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_14_n104), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_14_n107) );
  OAI211_X1 SD1_SB_inst_SD1_SB_bit_inst_14_U15 ( .C1(CipherErrorVec[24]), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_14_n105), .A(
        SD1_SB_inst_SD1_SB_bit_inst_14_n99), .B(
        SD1_SB_inst_SD1_SB_bit_inst_14_n102), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_14_n109) );
  NAND3_X1 SD1_SB_inst_SD1_SB_bit_inst_14_U14 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_14_n101), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_14_n105), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_14_n100), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_14_n128) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_14_U13 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_14_n106), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_14_n105) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_14_U12 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_14_n104), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_14_n103) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_14_U11 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_14_n102), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_14_n101) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_14_U10 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_14_n100), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_14_n99) );
  MUX2_X1 SD1_SB_inst_SD1_SB_bit_inst_14_U9 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_14_n97), .B(
        SD1_SB_inst_SD1_SB_bit_inst_14_n98), .S(
        SD1_SB_inst_SD1_SB_bit_inst_14_n99), .Z(
        SD1_SB_inst_SD1_SB_bit_inst_14_n125) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_14_U8 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_14_n118), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_14_n97) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_14_U7 ( .A(CipherErrorVec[25]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_14_n104) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_14_U6 ( .A(CipherErrorVec[23]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_14_n102) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_14_U5 ( .A(CipherErrorVec[26]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_14_n106) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_14_U4 ( .A(CipherErrorVec[22]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_14_n100) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_14_U3 ( .A1(CipherErrorVec[24]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_14_n121), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_14_n98) );
  AOI222_X1 SD1_SB_inst_SD1_SB_bit_inst_15_U45 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_15_n141), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_15_n140), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_15_n141), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_15_n139), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_15_n140), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_15_n138), .ZN(Feedback[59]) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_15_U44 ( .A(StateRegOutput[12]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_15_n137), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_15_n138) );
  AOI211_X1 SD1_SB_inst_SD1_SB_bit_inst_15_U43 ( .C1(
        SD1_SB_inst_SD1_SB_bit_inst_15_n136), .C2(CipherErrorVec[24]), .A(
        SD1_SB_inst_SD1_SB_bit_inst_15_n135), .B(
        SD1_SB_inst_SD1_SB_bit_inst_15_n134), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_15_n137) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_15_U42 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_15_n105), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_15_n103), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_15_n133), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_15_n134) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_15_U41 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_15_n107), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_15_n132), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_15_n131), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_15_n135) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_15_U40 ( .A1(CipherErrorVec[24]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_15_n100), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_15_n131) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_15_U39 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_15_n130), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_15_n136) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_15_U38 ( .A(StateRegOutput[14]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_15_n129), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_15_n139) );
  AOI22_X1 SD1_SB_inst_SD1_SB_bit_inst_15_U37 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_15_n128), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_15_n127), .B1(CipherErrorVec[27]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_15_n126), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_15_n129) );
  OAI211_X1 SD1_SB_inst_SD1_SB_bit_inst_15_U36 ( .C1(
        SD1_SB_inst_SD1_SB_bit_inst_15_n125), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_15_n101), .A(
        SD1_SB_inst_SD1_SB_bit_inst_15_n124), .B(
        SD1_SB_inst_SD1_SB_bit_inst_15_n123), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_15_n126) );
  NAND3_X1 SD1_SB_inst_SD1_SB_bit_inst_15_U35 ( .A1(CipherErrorVec[21]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_15_n108), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_15_n122), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_15_n123) );
  OAI22_X1 SD1_SB_inst_SD1_SB_bit_inst_15_U34 ( .A1(CipherErrorVec[24]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_15_n106), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_15_n100), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_15_n103), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_15_n122) );
  AOI22_X1 SD1_SB_inst_SD1_SB_bit_inst_15_U33 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_15_n102), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_15_n104), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_15_n105), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_15_n108), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_15_n125) );
  OAI21_X1 SD1_SB_inst_SD1_SB_bit_inst_15_U32 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_15_n100), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_15_n121), .A(
        SD1_SB_inst_SD1_SB_bit_inst_15_n120), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_15_n127) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_15_U31 ( .A(CipherErrorVec[21]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_15_n121) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_15_U30 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_15_n124), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_15_n128) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_15_U29 ( .A(StateRegOutput[13]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_15_n119), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_15_n140) );
  AOI22_X1 SD1_SB_inst_SD1_SB_bit_inst_15_U28 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_15_n105), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_15_n118), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_15_n100), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_15_n117), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_15_n119) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_15_U27 ( .A1(CipherErrorVec[24]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_15_n132), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_15_n108), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_15_n117) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_15_U26 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_15_n102), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_15_n105), .A3(CipherErrorVec[21]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_15_n132) );
  OAI22_X1 SD1_SB_inst_SD1_SB_bit_inst_15_U25 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_15_n102), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_15_n133), .B1(CipherErrorVec[27]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_15_n130), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_15_n118) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_15_U24 ( .A1(CipherErrorVec[21]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_15_n116), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_15_n133) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_15_U23 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_15_n115), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_15_n101), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_15_n116) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_15_U22 ( .A1(CipherErrorVec[24]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_15_n107), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_15_n115) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_15_U21 ( .A(StateRegOutput[15]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_15_n114), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_15_n141) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_15_U20 ( .B1(CipherErrorVec[27]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_15_n113), .A(
        SD1_SB_inst_SD1_SB_bit_inst_15_n112), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_15_n114) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_15_U19 ( .B1(CipherErrorVec[21]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_15_n124), .A(
        SD1_SB_inst_SD1_SB_bit_inst_15_n120), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_15_n112) );
  NAND3_X1 SD1_SB_inst_SD1_SB_bit_inst_15_U18 ( .A1(CipherErrorVec[24]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_15_n100), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_15_n107), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_15_n120) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_15_U17 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_15_n102), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_15_n105), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_15_n124) );
  OAI221_X1 SD1_SB_inst_SD1_SB_bit_inst_15_U16 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_15_n105), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_15_n130), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_15_n105), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_15_n111), .A(
        SD1_SB_inst_SD1_SB_bit_inst_15_n110), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_15_n113) );
  OAI21_X1 SD1_SB_inst_SD1_SB_bit_inst_15_U15 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_15_n107), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_15_n109), .A(CipherErrorVec[24]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_15_n110) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_15_U14 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_15_n102), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_15_n100), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_15_n106), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_15_n109) );
  OAI211_X1 SD1_SB_inst_SD1_SB_bit_inst_15_U13 ( .C1(CipherErrorVec[24]), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_15_n107), .A(
        SD1_SB_inst_SD1_SB_bit_inst_15_n100), .B(
        SD1_SB_inst_SD1_SB_bit_inst_15_n103), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_15_n111) );
  NAND3_X1 SD1_SB_inst_SD1_SB_bit_inst_15_U12 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_15_n102), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_15_n107), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_15_n101), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_15_n130) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_15_U11 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_15_n108), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_15_n107) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_15_U10 ( .A(CipherErrorVec[25]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_15_n106) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_15_U9 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_15_n106), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_15_n105) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_15_U8 ( .A(CipherErrorVec[24]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_15_n104) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_15_U7 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_15_n103), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_15_n102) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_15_U6 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_15_n101), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_15_n100) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_15_U5 ( .A(CipherErrorVec[23]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_15_n103) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_15_U4 ( .A(CipherErrorVec[26]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_15_n108) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_15_U3 ( .A(CipherErrorVec[22]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_15_n101) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_16_U48 ( .B1(OutputRegIn[18]), .B2(
        OutputRegIn[19]), .A(SD1_SB_inst_SD1_SB_bit_inst_16_n132), .ZN(
        Feedback[32]) );
  AOI221_X1 SD1_SB_inst_SD1_SB_bit_inst_16_U47 ( .B1(OutputRegIn[18]), .B2(
        OutputRegIn[16]), .C1(OutputRegIn[19]), .C2(OutputRegIn[16]), .A(
        OutputRegIn[17]), .ZN(SD1_SB_inst_SD1_SB_bit_inst_16_n132) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_16_U46 ( .A(StateRegOutput[17]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_16_n131), .ZN(OutputRegIn[17]) );
  AOI221_X1 SD1_SB_inst_SD1_SB_bit_inst_16_U45 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_16_n130), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_16_n104), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_16_n129), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_16_n104), .A(
        SD1_SB_inst_SD1_SB_bit_inst_16_n128), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_16_n131) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_16_U44 ( .A1(CipherErrorVec[30]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_16_n103), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_16_n127), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_16_n128) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_16_U43 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_16_n100), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_16_n126), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_16_n129) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_16_U42 ( .A1(CipherErrorVec[34]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_16_n125), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_16_n130) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_16_U41 ( .A(StateRegOutput[19]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_16_n124), .ZN(OutputRegIn[19]) );
  AOI211_X1 SD1_SB_inst_SD1_SB_bit_inst_16_U40 ( .C1(CipherErrorVec[34]), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_16_n123), .A(
        SD1_SB_inst_SD1_SB_bit_inst_16_n122), .B(
        SD1_SB_inst_SD1_SB_bit_inst_16_n121), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_16_n124) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_16_U39 ( .A1(CipherErrorVec[28]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_16_n98), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_16_n120), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_16_n121) );
  AOI222_X1 SD1_SB_inst_SD1_SB_bit_inst_16_U38 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_16_n105), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_16_n101), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_16_n105), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_16_n119), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_16_n101), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_16_n118), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_16_n123) );
  OAI221_X1 SD1_SB_inst_SD1_SB_bit_inst_16_U37 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_16_n117), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_16_n97), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_16_n117), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_16_n99), .A(
        SD1_SB_inst_SD1_SB_bit_inst_16_n103), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_16_n118) );
  OAI211_X1 SD1_SB_inst_SD1_SB_bit_inst_16_U36 ( .C1(
        SD1_SB_inst_SD1_SB_bit_inst_16_n102), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_16_n97), .A(
        SD1_SB_inst_SD1_SB_bit_inst_16_n116), .B(
        SD1_SB_inst_SD1_SB_bit_inst_16_n99), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_16_n119) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_16_U35 ( .A(StateRegOutput[18]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_16_n115), .ZN(OutputRegIn[18]) );
  AOI211_X1 SD1_SB_inst_SD1_SB_bit_inst_16_U34 ( .C1(CipherErrorVec[34]), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_16_n114), .A(
        SD1_SB_inst_SD1_SB_bit_inst_16_n122), .B(
        SD1_SB_inst_SD1_SB_bit_inst_16_n113), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_16_n115) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_16_U33 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_16_n125), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_16_n93), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_16_n113) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_16_U32 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_16_n102), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_16_n117), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_16_n125) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_16_U31 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_16_n99), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_16_n120), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_16_n116), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_16_n122) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_16_U30 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_16_n102), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_16_n97), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_16_n116) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_16_U29 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_16_n104), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_16_n100), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_16_n120) );
  OAI22_X1 SD1_SB_inst_SD1_SB_bit_inst_16_U28 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_16_n104), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_16_n112), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_16_n111), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_16_n99), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_16_n114) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_16_U27 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_16_n97), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_16_n101), .A(
        SD1_SB_inst_SD1_SB_bit_inst_16_n102), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_16_n111) );
  AOI22_X1 SD1_SB_inst_SD1_SB_bit_inst_16_U26 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_16_n102), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_16_n97), .B1(CipherErrorVec[28]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_16_n110), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_16_n112) );
  OAI21_X1 SD1_SB_inst_SD1_SB_bit_inst_16_U25 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_16_n100), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_16_n103), .A(
        SD1_SB_inst_SD1_SB_bit_inst_16_n109), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_16_n110) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_16_U24 ( .A(StateRegOutput[16]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_16_n108), .ZN(OutputRegIn[16]) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_16_U23 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_16_n107), .B2(CipherErrorVec[30]), .A(
        SD1_SB_inst_SD1_SB_bit_inst_16_n106), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_16_n108) );
  AOI221_X1 SD1_SB_inst_SD1_SB_bit_inst_16_U22 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_16_n104), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_16_n109), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_16_n105), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_16_n126), .A(
        SD1_SB_inst_SD1_SB_bit_inst_16_n101), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_16_n106) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_16_U21 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_16_n117), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_16_n109) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_16_U20 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_16_n97), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_16_n99), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_16_n117) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_16_U19 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_16_n127), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_16_n102), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_16_n107) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_16_U18 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_16_n105), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_16_n104) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_16_U17 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_16_n103), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_16_n102) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_16_U16 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_16_n101), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_16_n100) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_16_U15 ( .A(CipherErrorVec[30]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_16_n99) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_16_U14 ( .A(CipherErrorVec[29]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_16_n98) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_16_U13 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_16_n98), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_16_n97) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_16_U12 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_16_n96), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_16_n127) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_16_U11 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_16_n94), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_16_n126) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_16_U10 ( .A(CipherErrorVec[28]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_16_n93) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_16_U9 ( .A(CipherErrorVec[33]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_16_n105) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_16_U8 ( .A(CipherErrorVec[32]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_16_n103) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_16_U7 ( .A(CipherErrorVec[31]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_16_n101) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_16_U6 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_16_n97), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_16_n104), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_16_n95) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_16_U5 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_16_n95), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_16_n101), .A(
        SD1_SB_inst_SD1_SB_bit_inst_16_n93), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_16_n96) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_16_U4 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_16_n102), .A2(CipherErrorVec[30]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_16_n92) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_16_U3 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_16_n92), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_16_n93), .A(
        SD1_SB_inst_SD1_SB_bit_inst_16_n98), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_16_n94) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_17_U36 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_17_n109), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_17_n108), .A(
        SD1_SB_inst_SD1_SB_bit_inst_17_n107), .ZN(Feedback[33]) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_17_U35 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_17_n106), .B2(StateRegOutput[16]), .A(
        SD1_SB_inst_SD1_SB_bit_inst_17_n105), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_17_n107) );
  OAI22_X1 SD1_SB_inst_SD1_SB_bit_inst_17_U34 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_17_n108), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_17_n109), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_17_n106), .B2(StateRegOutput[16]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_17_n105) );
  AOI22_X1 SD1_SB_inst_SD1_SB_bit_inst_17_U33 ( .A1(CipherErrorVec[28]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_17_n104), .B1(CipherErrorVec[31]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_17_n103), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_17_n106) );
  OAI21_X1 SD1_SB_inst_SD1_SB_bit_inst_17_U32 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_17_n102), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_17_n101), .A(
        SD1_SB_inst_SD1_SB_bit_inst_17_n100), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_17_n103) );
  NAND3_X1 SD1_SB_inst_SD1_SB_bit_inst_17_U31 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_17_n86), .A2(CipherErrorVec[33]), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_17_n85), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_17_n100) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_17_U30 ( .A1(CipherErrorVec[28]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_17_n86), .A3(CipherErrorVec[32]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_17_n102) );
  AOI211_X1 SD1_SB_inst_SD1_SB_bit_inst_17_U29 ( .C1(
        SD1_SB_inst_SD1_SB_bit_inst_17_n99), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_17_n85), .A(CipherErrorVec[32]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_17_n87), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_17_n104) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_17_U28 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_17_n84), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_17_n90), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_17_n101) );
  XOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_17_U27 ( .A(StateRegOutput[19]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_17_n95), .Z(
        SD1_SB_inst_SD1_SB_bit_inst_17_n109) );
  OAI21_X1 SD1_SB_inst_SD1_SB_bit_inst_17_U26 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_17_n94), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_17_n98), .A(
        SD1_SB_inst_SD1_SB_bit_inst_17_n93), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_17_n95) );
  OAI221_X1 SD1_SB_inst_SD1_SB_bit_inst_17_U25 ( .B1(CipherErrorVec[32]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_17_n92), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_17_n89), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_17_n91), .A(CipherErrorVec[34]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_17_n93) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_17_U24 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_17_n84), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_17_n86), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_17_n88), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_17_n91) );
  OAI33_X1 SD1_SB_inst_SD1_SB_bit_inst_17_U23 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_17_n86), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_17_n99), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_17_n85), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_17_n87), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_17_n90), .B3(
        SD1_SB_inst_SD1_SB_bit_inst_17_n84), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_17_n92) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_17_U22 ( .A1(CipherErrorVec[31]), .A2(
        CipherErrorVec[33]), .ZN(SD1_SB_inst_SD1_SB_bit_inst_17_n99) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_17_U21 ( .A1(CipherErrorVec[31]), .A2(
        CipherErrorVec[33]), .ZN(SD1_SB_inst_SD1_SB_bit_inst_17_n98) );
  AOI221_X1 SD1_SB_inst_SD1_SB_bit_inst_17_U20 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_17_n96), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_17_n84), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_17_n97), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_17_n84), .A(CipherErrorVec[34]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_17_n94) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_17_U19 ( .A(CipherErrorVec[28]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_17_n97) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_17_U18 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_17_n87), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_17_n89), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_17_n96) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_17_U17 ( .A(CipherErrorVec[31]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_17_n88) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_17_U16 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_17_n87), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_17_n86) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_17_U15 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_17_n85), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_17_n84) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_17_U14 ( .A(CipherErrorVec[32]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_17_n89) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_17_U13 ( .A(CipherErrorVec[33]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_17_n90) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_17_U12 ( .A(CipherErrorVec[30]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_17_n87) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_17_U11 ( .A(CipherErrorVec[29]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_17_n85) );
  XOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_17_U10 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_17_n83), .B(StateRegOutput[18]), .Z(
        SD1_SB_inst_SD1_SB_bit_inst_17_n108) );
  AOI22_X1 SD1_SB_inst_SD1_SB_bit_inst_17_U9 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_17_n77), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_17_n96), .B1(CipherErrorVec[34]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_17_n82), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_17_n83) );
  OAI22_X1 SD1_SB_inst_SD1_SB_bit_inst_17_U8 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_17_n87), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_17_n79), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_17_n89), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_17_n81), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_17_n82) );
  AOI211_X1 SD1_SB_inst_SD1_SB_bit_inst_17_U7 ( .C1(CipherErrorVec[28]), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_17_n99), .A(
        SD1_SB_inst_SD1_SB_bit_inst_17_n86), .B(
        SD1_SB_inst_SD1_SB_bit_inst_17_n80), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_17_n81) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_17_U6 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_17_n101), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_17_n80) );
  AOI22_X1 SD1_SB_inst_SD1_SB_bit_inst_17_U5 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_17_n84), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_17_n88), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_17_n90), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_17_n78), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_17_n79) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_17_U4 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_17_n84), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_17_n97), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_17_n78) );
  AOI22_X1 SD1_SB_inst_SD1_SB_bit_inst_17_U3 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_17_n84), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_17_n98), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_17_n85), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_17_n97), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_17_n77) );
  OAI22_X1 SD1_SB_inst_SD1_SB_bit_inst_18_U44 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_18_n137), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_18_n136), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_18_n135), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_18_n134), .ZN(Feedback[34]) );
  XOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_18_U43 ( .A(StateRegOutput[17]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_18_n133), .Z(
        SD1_SB_inst_SD1_SB_bit_inst_18_n136) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_18_U42 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_18_n110), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_18_n132), .A(
        SD1_SB_inst_SD1_SB_bit_inst_18_n131), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_18_n133) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_18_U41 ( .A1(CipherErrorVec[31]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_18_n130), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_18_n129), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_18_n131) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_18_U40 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_18_n112), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_18_n106), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_18_n129) );
  OAI22_X1 SD1_SB_inst_SD1_SB_bit_inst_18_U39 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_18_n108), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_18_n128), .B1(CipherErrorVec[34]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_18_n127), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_18_n132) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_18_U38 ( .A(StateRegOutput[16]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_18_n124), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_18_n135) );
  AOI22_X1 SD1_SB_inst_SD1_SB_bit_inst_18_U37 ( .A1(CipherErrorVec[31]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_18_n123), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_18_n108), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_18_n122), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_18_n124) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_18_U36 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_18_n110), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_18_n128), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_18_n122) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_18_U35 ( .A1(CipherErrorVec[28]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_18_n121), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_18_n128) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_18_U34 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_18_n126), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_18_n107), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_18_n121) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_18_U33 ( .A1(CipherErrorVec[31]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_18_n112), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_18_n126) );
  OAI21_X1 SD1_SB_inst_SD1_SB_bit_inst_18_U32 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_18_n130), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_18_n120), .A(
        SD1_SB_inst_SD1_SB_bit_inst_18_n127), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_18_n123) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_18_U31 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_18_n106), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_18_n113), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_18_n120) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_18_U30 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_18_n108), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_18_n110), .A3(CipherErrorVec[28]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_18_n130) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_18_U29 ( .A(StateRegOutput[19]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_18_n119), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_18_n134) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_18_U28 ( .B1(CipherErrorVec[34]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_18_n118), .A(
        SD1_SB_inst_SD1_SB_bit_inst_18_n117), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_18_n119) );
  AOI221_X1 SD1_SB_inst_SD1_SB_bit_inst_18_U27 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_18_n111), .B2(CipherErrorVec[28]), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_18_n109), .C2(CipherErrorVec[28]), .A(
        SD1_SB_inst_SD1_SB_bit_inst_18_n125), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_18_n117) );
  NAND3_X1 SD1_SB_inst_SD1_SB_bit_inst_18_U26 ( .A1(CipherErrorVec[31]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_18_n112), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_18_n106), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_18_n125) );
  OAI221_X1 SD1_SB_inst_SD1_SB_bit_inst_18_U25 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_18_n110), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_18_n127), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_18_n110), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_18_n116), .A(
        SD1_SB_inst_SD1_SB_bit_inst_18_n115), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_18_n118) );
  OAI21_X1 SD1_SB_inst_SD1_SB_bit_inst_18_U24 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_18_n112), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_18_n114), .A(CipherErrorVec[31]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_18_n115) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_18_U23 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_18_n108), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_18_n106), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_18_n111), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_18_n114) );
  OAI211_X1 SD1_SB_inst_SD1_SB_bit_inst_18_U22 ( .C1(CipherErrorVec[31]), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_18_n112), .A(
        SD1_SB_inst_SD1_SB_bit_inst_18_n106), .B(
        SD1_SB_inst_SD1_SB_bit_inst_18_n109), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_18_n116) );
  NAND3_X1 SD1_SB_inst_SD1_SB_bit_inst_18_U21 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_18_n108), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_18_n112), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_18_n107), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_18_n127) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_18_U20 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_18_n113), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_18_n112) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_18_U19 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_18_n111), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_18_n110) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_18_U18 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_18_n109), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_18_n108) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_18_U17 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_18_n107), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_18_n106) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_18_U16 ( .A(CipherErrorVec[32]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_18_n111) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_18_U15 ( .A(CipherErrorVec[30]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_18_n109) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_18_U14 ( .A(CipherErrorVec[33]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_18_n113) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_18_U13 ( .A(CipherErrorVec[29]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_18_n107) );
  AOI221_X1 SD1_SB_inst_SD1_SB_bit_inst_18_U12 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_18_n135), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_18_n134), .C1(StateRegOutput[18]), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_18_n104), .A(
        SD1_SB_inst_SD1_SB_bit_inst_18_n105), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_18_n137) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_18_U11 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_18_n104), .A2(StateRegOutput[18]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_18_n105) );
  AOI211_X1 SD1_SB_inst_SD1_SB_bit_inst_18_U10 ( .C1(
        SD1_SB_inst_SD1_SB_bit_inst_18_n108), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_18_n99), .A(
        SD1_SB_inst_SD1_SB_bit_inst_18_n102), .B(
        SD1_SB_inst_SD1_SB_bit_inst_18_n103), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_18_n104) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_18_U9 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_18_n111), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_18_n109), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_18_n125), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_18_n103) );
  AOI211_X1 SD1_SB_inst_SD1_SB_bit_inst_18_U8 ( .C1(
        SD1_SB_inst_SD1_SB_bit_inst_18_n109), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_18_n100), .A(
        SD1_SB_inst_SD1_SB_bit_inst_18_n111), .B(
        SD1_SB_inst_SD1_SB_bit_inst_18_n101), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_18_n102) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_18_U7 ( .A(CipherErrorVec[34]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_18_n101) );
  AOI22_X1 SD1_SB_inst_SD1_SB_bit_inst_18_U6 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_18_n106), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_18_n113), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_18_n126), .B2(CipherErrorVec[28]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_18_n100) );
  OAI22_X1 SD1_SB_inst_SD1_SB_bit_inst_18_U5 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_18_n106), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_18_n97), .B1(CipherErrorVec[31]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_18_n98), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_18_n99) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_18_U4 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_18_n106), .A2(CipherErrorVec[34]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_18_n98) );
  OAI221_X1 SD1_SB_inst_SD1_SB_bit_inst_18_U3 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_18_n110), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_18_n113), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_18_n110), .C2(CipherErrorVec[34]), .A(
        CipherErrorVec[28]), .ZN(SD1_SB_inst_SD1_SB_bit_inst_18_n97) );
  AOI222_X1 SD1_SB_inst_SD1_SB_bit_inst_19_U45 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_19_n141), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_19_n140), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_19_n141), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_19_n139), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_19_n140), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_19_n138), .ZN(Feedback[35]) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_19_U44 ( .A(StateRegOutput[16]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_19_n137), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_19_n138) );
  AOI211_X1 SD1_SB_inst_SD1_SB_bit_inst_19_U43 ( .C1(
        SD1_SB_inst_SD1_SB_bit_inst_19_n136), .C2(CipherErrorVec[31]), .A(
        SD1_SB_inst_SD1_SB_bit_inst_19_n135), .B(
        SD1_SB_inst_SD1_SB_bit_inst_19_n134), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_19_n137) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_19_U42 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_19_n105), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_19_n103), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_19_n133), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_19_n134) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_19_U41 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_19_n107), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_19_n132), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_19_n131), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_19_n135) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_19_U40 ( .A1(CipherErrorVec[31]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_19_n100), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_19_n131) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_19_U39 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_19_n130), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_19_n136) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_19_U38 ( .A(StateRegOutput[18]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_19_n129), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_19_n139) );
  AOI22_X1 SD1_SB_inst_SD1_SB_bit_inst_19_U37 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_19_n128), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_19_n127), .B1(CipherErrorVec[34]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_19_n126), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_19_n129) );
  OAI211_X1 SD1_SB_inst_SD1_SB_bit_inst_19_U36 ( .C1(
        SD1_SB_inst_SD1_SB_bit_inst_19_n125), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_19_n101), .A(
        SD1_SB_inst_SD1_SB_bit_inst_19_n124), .B(
        SD1_SB_inst_SD1_SB_bit_inst_19_n123), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_19_n126) );
  NAND3_X1 SD1_SB_inst_SD1_SB_bit_inst_19_U35 ( .A1(CipherErrorVec[28]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_19_n108), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_19_n122), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_19_n123) );
  OAI22_X1 SD1_SB_inst_SD1_SB_bit_inst_19_U34 ( .A1(CipherErrorVec[31]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_19_n106), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_19_n100), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_19_n103), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_19_n122) );
  AOI22_X1 SD1_SB_inst_SD1_SB_bit_inst_19_U33 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_19_n102), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_19_n104), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_19_n105), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_19_n108), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_19_n125) );
  OAI21_X1 SD1_SB_inst_SD1_SB_bit_inst_19_U32 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_19_n100), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_19_n121), .A(
        SD1_SB_inst_SD1_SB_bit_inst_19_n120), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_19_n127) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_19_U31 ( .A(CipherErrorVec[28]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_19_n121) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_19_U30 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_19_n124), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_19_n128) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_19_U29 ( .A(StateRegOutput[17]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_19_n119), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_19_n140) );
  AOI22_X1 SD1_SB_inst_SD1_SB_bit_inst_19_U28 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_19_n105), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_19_n118), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_19_n100), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_19_n117), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_19_n119) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_19_U27 ( .A1(CipherErrorVec[31]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_19_n132), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_19_n108), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_19_n117) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_19_U26 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_19_n102), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_19_n105), .A3(CipherErrorVec[28]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_19_n132) );
  OAI22_X1 SD1_SB_inst_SD1_SB_bit_inst_19_U25 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_19_n102), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_19_n133), .B1(CipherErrorVec[34]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_19_n130), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_19_n118) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_19_U24 ( .A1(CipherErrorVec[28]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_19_n116), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_19_n133) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_19_U23 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_19_n115), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_19_n101), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_19_n116) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_19_U22 ( .A1(CipherErrorVec[31]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_19_n107), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_19_n115) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_19_U21 ( .A(StateRegOutput[19]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_19_n114), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_19_n141) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_19_U20 ( .B1(CipherErrorVec[34]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_19_n113), .A(
        SD1_SB_inst_SD1_SB_bit_inst_19_n112), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_19_n114) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_19_U19 ( .B1(CipherErrorVec[28]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_19_n124), .A(
        SD1_SB_inst_SD1_SB_bit_inst_19_n120), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_19_n112) );
  NAND3_X1 SD1_SB_inst_SD1_SB_bit_inst_19_U18 ( .A1(CipherErrorVec[31]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_19_n100), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_19_n107), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_19_n120) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_19_U17 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_19_n102), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_19_n105), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_19_n124) );
  OAI221_X1 SD1_SB_inst_SD1_SB_bit_inst_19_U16 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_19_n105), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_19_n130), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_19_n105), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_19_n111), .A(
        SD1_SB_inst_SD1_SB_bit_inst_19_n110), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_19_n113) );
  OAI21_X1 SD1_SB_inst_SD1_SB_bit_inst_19_U15 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_19_n107), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_19_n109), .A(CipherErrorVec[31]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_19_n110) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_19_U14 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_19_n102), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_19_n100), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_19_n106), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_19_n109) );
  OAI211_X1 SD1_SB_inst_SD1_SB_bit_inst_19_U13 ( .C1(CipherErrorVec[31]), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_19_n107), .A(
        SD1_SB_inst_SD1_SB_bit_inst_19_n100), .B(
        SD1_SB_inst_SD1_SB_bit_inst_19_n103), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_19_n111) );
  NAND3_X1 SD1_SB_inst_SD1_SB_bit_inst_19_U12 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_19_n102), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_19_n107), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_19_n101), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_19_n130) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_19_U11 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_19_n108), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_19_n107) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_19_U10 ( .A(CipherErrorVec[32]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_19_n106) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_19_U9 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_19_n106), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_19_n105) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_19_U8 ( .A(CipherErrorVec[31]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_19_n104) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_19_U7 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_19_n103), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_19_n102) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_19_U6 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_19_n101), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_19_n100) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_19_U5 ( .A(CipherErrorVec[30]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_19_n103) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_19_U4 ( .A(CipherErrorVec[33]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_19_n108) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_19_U3 ( .A(CipherErrorVec[29]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_19_n101) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_20_U47 ( .B1(OutputRegIn[22]), .B2(
        OutputRegIn[23]), .A(SD1_SB_inst_SD1_SB_bit_inst_20_n131), .ZN(
        Feedback[44]) );
  AOI221_X1 SD1_SB_inst_SD1_SB_bit_inst_20_U46 ( .B1(OutputRegIn[22]), .B2(
        OutputRegIn[20]), .C1(OutputRegIn[23]), .C2(OutputRegIn[20]), .A(
        OutputRegIn[21]), .ZN(SD1_SB_inst_SD1_SB_bit_inst_20_n131) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_20_U45 ( .A(StateRegOutput[23]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_20_n127), .ZN(OutputRegIn[23]) );
  AOI211_X1 SD1_SB_inst_SD1_SB_bit_inst_20_U44 ( .C1(CipherErrorVec[41]), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_20_n126), .A(
        SD1_SB_inst_SD1_SB_bit_inst_20_n125), .B(
        SD1_SB_inst_SD1_SB_bit_inst_20_n124), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_20_n127) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_20_U43 ( .A1(CipherErrorVec[35]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_20_n101), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_20_n123), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_20_n124) );
  AOI222_X1 SD1_SB_inst_SD1_SB_bit_inst_20_U42 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_20_n108), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_20_n104), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_20_n108), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_20_n122), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_20_n104), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_20_n121), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_20_n126) );
  OAI221_X1 SD1_SB_inst_SD1_SB_bit_inst_20_U41 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_20_n120), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_20_n100), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_20_n120), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_20_n102), .A(
        SD1_SB_inst_SD1_SB_bit_inst_20_n106), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_20_n121) );
  OAI211_X1 SD1_SB_inst_SD1_SB_bit_inst_20_U40 ( .C1(
        SD1_SB_inst_SD1_SB_bit_inst_20_n105), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_20_n100), .A(
        SD1_SB_inst_SD1_SB_bit_inst_20_n119), .B(
        SD1_SB_inst_SD1_SB_bit_inst_20_n102), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_20_n122) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_20_U39 ( .A(StateRegOutput[22]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_20_n118), .ZN(OutputRegIn[22]) );
  AOI211_X1 SD1_SB_inst_SD1_SB_bit_inst_20_U38 ( .C1(CipherErrorVec[41]), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_20_n117), .A(
        SD1_SB_inst_SD1_SB_bit_inst_20_n125), .B(
        SD1_SB_inst_SD1_SB_bit_inst_20_n116), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_20_n118) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_20_U37 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_20_n128), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_20_n96), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_20_n116) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_20_U36 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_20_n105), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_20_n120), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_20_n128) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_20_U35 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_20_n102), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_20_n123), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_20_n119), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_20_n125) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_20_U34 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_20_n105), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_20_n100), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_20_n119) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_20_U33 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_20_n107), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_20_n103), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_20_n123) );
  OAI22_X1 SD1_SB_inst_SD1_SB_bit_inst_20_U32 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_20_n107), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_20_n115), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_20_n114), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_20_n102), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_20_n117) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_20_U31 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_20_n100), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_20_n104), .A(
        SD1_SB_inst_SD1_SB_bit_inst_20_n105), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_20_n114) );
  AOI22_X1 SD1_SB_inst_SD1_SB_bit_inst_20_U30 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_20_n105), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_20_n100), .B1(CipherErrorVec[35]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_20_n113), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_20_n115) );
  OAI21_X1 SD1_SB_inst_SD1_SB_bit_inst_20_U29 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_20_n103), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_20_n106), .A(
        SD1_SB_inst_SD1_SB_bit_inst_20_n112), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_20_n113) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_20_U28 ( .A(StateRegOutput[20]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_20_n111), .ZN(OutputRegIn[20]) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_20_U27 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_20_n110), .B2(CipherErrorVec[37]), .A(
        SD1_SB_inst_SD1_SB_bit_inst_20_n109), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_20_n111) );
  AOI221_X1 SD1_SB_inst_SD1_SB_bit_inst_20_U26 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_20_n107), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_20_n112), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_20_n108), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_20_n129), .A(
        SD1_SB_inst_SD1_SB_bit_inst_20_n104), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_20_n109) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_20_U25 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_20_n120), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_20_n112) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_20_U24 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_20_n100), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_20_n102), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_20_n120) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_20_U23 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_20_n130), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_20_n105), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_20_n110) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_20_U22 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_20_n108), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_20_n107) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_20_U21 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_20_n106), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_20_n105) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_20_U20 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_20_n104), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_20_n103) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_20_U19 ( .A(CipherErrorVec[37]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_20_n102) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_20_U18 ( .A(CipherErrorVec[36]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_20_n101) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_20_U17 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_20_n101), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_20_n100) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_20_U16 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_20_n99), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_20_n130) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_20_U15 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_20_n97), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_20_n129) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_20_U14 ( .A(CipherErrorVec[35]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_20_n96) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_20_U13 ( .A(CipherErrorVec[40]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_20_n108) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_20_U12 ( .A(CipherErrorVec[39]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_20_n106) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_20_U11 ( .A(CipherErrorVec[38]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_20_n104) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_20_U10 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_20_n100), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_20_n107), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_20_n98) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_20_U9 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_20_n98), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_20_n104), .A(
        SD1_SB_inst_SD1_SB_bit_inst_20_n96), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_20_n99) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_20_U8 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_20_n105), .A2(CipherErrorVec[37]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_20_n95) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_20_U7 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_20_n95), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_20_n96), .A(
        SD1_SB_inst_SD1_SB_bit_inst_20_n101), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_20_n97) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_20_U6 ( .A(StateRegOutput[21]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_20_n94), .ZN(OutputRegIn[21]) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_20_U5 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_20_n107), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_20_n92), .A(
        SD1_SB_inst_SD1_SB_bit_inst_20_n93), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_20_n94) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_20_U4 ( .A1(CipherErrorVec[37]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_20_n130), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_20_n106), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_20_n93) );
  OAI22_X1 SD1_SB_inst_SD1_SB_bit_inst_20_U3 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_20_n103), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_20_n129), .B1(CipherErrorVec[41]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_20_n128), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_20_n92) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_21_U37 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_21_n110), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_21_n109), .A(
        SD1_SB_inst_SD1_SB_bit_inst_21_n108), .ZN(Feedback[45]) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_21_U36 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_21_n107), .B2(StateRegOutput[20]), .A(
        SD1_SB_inst_SD1_SB_bit_inst_21_n106), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_21_n108) );
  OAI22_X1 SD1_SB_inst_SD1_SB_bit_inst_21_U35 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_21_n109), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_21_n110), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_21_n107), .B2(StateRegOutput[20]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_21_n106) );
  AOI22_X1 SD1_SB_inst_SD1_SB_bit_inst_21_U34 ( .A1(CipherErrorVec[35]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_21_n105), .B1(CipherErrorVec[38]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_21_n104), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_21_n107) );
  OAI21_X1 SD1_SB_inst_SD1_SB_bit_inst_21_U33 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_21_n103), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_21_n102), .A(
        SD1_SB_inst_SD1_SB_bit_inst_21_n101), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_21_n104) );
  NAND3_X1 SD1_SB_inst_SD1_SB_bit_inst_21_U32 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_21_n79), .A2(CipherErrorVec[40]), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_21_n78), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_21_n101) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_21_U31 ( .A1(CipherErrorVec[35]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_21_n79), .A3(CipherErrorVec[39]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_21_n103) );
  AOI211_X1 SD1_SB_inst_SD1_SB_bit_inst_21_U30 ( .C1(
        SD1_SB_inst_SD1_SB_bit_inst_21_n100), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_21_n78), .A(CipherErrorVec[39]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_21_n80), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_21_n105) );
  XOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_21_U29 ( .A(StateRegOutput[22]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_21_n99), .Z(
        SD1_SB_inst_SD1_SB_bit_inst_21_n109) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_21_U28 ( .B1(CipherErrorVec[41]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_21_n98), .A(
        SD1_SB_inst_SD1_SB_bit_inst_21_n97), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_21_n99) );
  AOI221_X1 SD1_SB_inst_SD1_SB_bit_inst_21_U27 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_21_n77), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_21_n96), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_21_n78), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_21_n95), .A(
        SD1_SB_inst_SD1_SB_bit_inst_21_n94), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_21_n97) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_21_U26 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_21_n93), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_21_n94) );
  OAI22_X1 SD1_SB_inst_SD1_SB_bit_inst_21_U25 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_21_n92), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_21_n80), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_21_n91), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_21_n82), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_21_n98) );
  AOI211_X1 SD1_SB_inst_SD1_SB_bit_inst_21_U24 ( .C1(CipherErrorVec[35]), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_21_n100), .A(
        SD1_SB_inst_SD1_SB_bit_inst_21_n79), .B(
        SD1_SB_inst_SD1_SB_bit_inst_21_n90), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_21_n91) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_21_U23 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_21_n102), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_21_n90) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_21_U22 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_21_n77), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_21_n83), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_21_n102) );
  AOI22_X1 SD1_SB_inst_SD1_SB_bit_inst_21_U21 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_21_n77), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_21_n81), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_21_n89), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_21_n83), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_21_n92) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_21_U20 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_21_n77), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_21_n95), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_21_n89) );
  XOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_21_U19 ( .A(StateRegOutput[23]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_21_n88), .Z(
        SD1_SB_inst_SD1_SB_bit_inst_21_n110) );
  OAI21_X1 SD1_SB_inst_SD1_SB_bit_inst_21_U18 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_21_n87), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_21_n96), .A(
        SD1_SB_inst_SD1_SB_bit_inst_21_n86), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_21_n88) );
  OAI221_X1 SD1_SB_inst_SD1_SB_bit_inst_21_U17 ( .B1(CipherErrorVec[39]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_21_n85), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_21_n82), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_21_n84), .A(CipherErrorVec[41]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_21_n86) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_21_U16 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_21_n77), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_21_n79), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_21_n81), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_21_n84) );
  OAI33_X1 SD1_SB_inst_SD1_SB_bit_inst_21_U15 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_21_n79), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_21_n100), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_21_n78), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_21_n80), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_21_n83), .B3(
        SD1_SB_inst_SD1_SB_bit_inst_21_n77), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_21_n85) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_21_U14 ( .A1(CipherErrorVec[38]), .A2(
        CipherErrorVec[40]), .ZN(SD1_SB_inst_SD1_SB_bit_inst_21_n100) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_21_U13 ( .A1(CipherErrorVec[38]), .A2(
        CipherErrorVec[40]), .ZN(SD1_SB_inst_SD1_SB_bit_inst_21_n96) );
  AOI221_X1 SD1_SB_inst_SD1_SB_bit_inst_21_U12 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_21_n93), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_21_n77), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_21_n95), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_21_n77), .A(CipherErrorVec[41]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_21_n87) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_21_U11 ( .A(CipherErrorVec[35]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_21_n95) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_21_U10 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_21_n80), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_21_n82), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_21_n93) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_21_U9 ( .A(CipherErrorVec[38]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_21_n81) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_21_U8 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_21_n80), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_21_n79) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_21_U7 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_21_n78), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_21_n77) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_21_U6 ( .A(CipherErrorVec[39]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_21_n82) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_21_U5 ( .A(CipherErrorVec[40]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_21_n83) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_21_U4 ( .A(CipherErrorVec[37]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_21_n80) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_21_U3 ( .A(CipherErrorVec[36]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_21_n78) );
  OAI22_X1 SD1_SB_inst_SD1_SB_bit_inst_22_U45 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_22_n138), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_22_n137), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_22_n136), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_22_n135), .ZN(Feedback[46]) );
  XOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_22_U44 ( .A(StateRegOutput[21]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_22_n134), .Z(
        SD1_SB_inst_SD1_SB_bit_inst_22_n137) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_22_U43 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_22_n103), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_22_n133), .A(
        SD1_SB_inst_SD1_SB_bit_inst_22_n132), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_22_n134) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_22_U42 ( .A1(CipherErrorVec[38]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_22_n131), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_22_n130), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_22_n132) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_22_U41 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_22_n105), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_22_n99), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_22_n130) );
  OAI22_X1 SD1_SB_inst_SD1_SB_bit_inst_22_U40 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_22_n101), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_22_n129), .B1(CipherErrorVec[41]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_22_n128), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_22_n133) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_22_U39 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_22_n135), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_22_n136), .A(
        SD1_SB_inst_SD1_SB_bit_inst_22_n127), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_22_n138) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_22_U38 ( .A(StateRegOutput[22]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_22_n126), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_22_n127) );
  AOI211_X1 SD1_SB_inst_SD1_SB_bit_inst_22_U37 ( .C1(
        SD1_SB_inst_SD1_SB_bit_inst_22_n101), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_22_n125), .A(
        SD1_SB_inst_SD1_SB_bit_inst_22_n124), .B(
        SD1_SB_inst_SD1_SB_bit_inst_22_n123), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_22_n126) );
  AOI211_X1 SD1_SB_inst_SD1_SB_bit_inst_22_U36 ( .C1(
        SD1_SB_inst_SD1_SB_bit_inst_22_n122), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_22_n102), .A(
        SD1_SB_inst_SD1_SB_bit_inst_22_n121), .B(
        SD1_SB_inst_SD1_SB_bit_inst_22_n104), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_22_n123) );
  AOI22_X1 SD1_SB_inst_SD1_SB_bit_inst_22_U35 ( .A1(CipherErrorVec[35]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_22_n120), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_22_n99), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_22_n106), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_22_n122) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_22_U34 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_22_n102), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_22_n104), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_22_n119), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_22_n124) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_22_U33 ( .A(CipherErrorVec[41]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_22_n121) );
  OAI221_X1 SD1_SB_inst_SD1_SB_bit_inst_22_U32 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_22_n103), .B2(CipherErrorVec[41]), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_22_n103), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_22_n106), .A(CipherErrorVec[35]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_22_n118) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_22_U31 ( .A(StateRegOutput[20]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_22_n117), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_22_n136) );
  AOI22_X1 SD1_SB_inst_SD1_SB_bit_inst_22_U30 ( .A1(CipherErrorVec[38]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_22_n116), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_22_n101), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_22_n115), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_22_n117) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_22_U29 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_22_n103), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_22_n129), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_22_n115) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_22_U28 ( .A1(CipherErrorVec[35]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_22_n114), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_22_n129) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_22_U27 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_22_n120), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_22_n100), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_22_n114) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_22_U26 ( .A1(CipherErrorVec[38]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_22_n105), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_22_n120) );
  OAI21_X1 SD1_SB_inst_SD1_SB_bit_inst_22_U25 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_22_n131), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_22_n113), .A(
        SD1_SB_inst_SD1_SB_bit_inst_22_n128), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_22_n116) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_22_U24 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_22_n99), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_22_n106), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_22_n113) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_22_U23 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_22_n101), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_22_n103), .A3(CipherErrorVec[35]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_22_n131) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_22_U22 ( .A(StateRegOutput[23]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_22_n112), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_22_n135) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_22_U21 ( .B1(CipherErrorVec[41]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_22_n111), .A(
        SD1_SB_inst_SD1_SB_bit_inst_22_n110), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_22_n112) );
  AOI221_X1 SD1_SB_inst_SD1_SB_bit_inst_22_U20 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_22_n104), .B2(CipherErrorVec[35]), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_22_n102), .C2(CipherErrorVec[35]), .A(
        SD1_SB_inst_SD1_SB_bit_inst_22_n119), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_22_n110) );
  NAND3_X1 SD1_SB_inst_SD1_SB_bit_inst_22_U19 ( .A1(CipherErrorVec[38]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_22_n105), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_22_n99), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_22_n119) );
  OAI221_X1 SD1_SB_inst_SD1_SB_bit_inst_22_U18 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_22_n103), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_22_n128), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_22_n103), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_22_n109), .A(
        SD1_SB_inst_SD1_SB_bit_inst_22_n108), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_22_n111) );
  OAI21_X1 SD1_SB_inst_SD1_SB_bit_inst_22_U17 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_22_n105), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_22_n107), .A(CipherErrorVec[38]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_22_n108) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_22_U16 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_22_n101), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_22_n99), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_22_n104), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_22_n107) );
  OAI211_X1 SD1_SB_inst_SD1_SB_bit_inst_22_U15 ( .C1(CipherErrorVec[38]), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_22_n105), .A(
        SD1_SB_inst_SD1_SB_bit_inst_22_n99), .B(
        SD1_SB_inst_SD1_SB_bit_inst_22_n102), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_22_n109) );
  NAND3_X1 SD1_SB_inst_SD1_SB_bit_inst_22_U14 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_22_n101), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_22_n105), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_22_n100), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_22_n128) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_22_U13 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_22_n106), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_22_n105) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_22_U12 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_22_n104), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_22_n103) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_22_U11 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_22_n102), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_22_n101) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_22_U10 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_22_n100), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_22_n99) );
  MUX2_X1 SD1_SB_inst_SD1_SB_bit_inst_22_U9 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_22_n97), .B(
        SD1_SB_inst_SD1_SB_bit_inst_22_n98), .S(
        SD1_SB_inst_SD1_SB_bit_inst_22_n99), .Z(
        SD1_SB_inst_SD1_SB_bit_inst_22_n125) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_22_U8 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_22_n118), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_22_n97) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_22_U7 ( .A(CipherErrorVec[39]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_22_n104) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_22_U6 ( .A(CipherErrorVec[37]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_22_n102) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_22_U5 ( .A(CipherErrorVec[40]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_22_n106) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_22_U4 ( .A(CipherErrorVec[36]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_22_n100) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_22_U3 ( .A1(CipherErrorVec[38]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_22_n121), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_22_n98) );
  AOI222_X1 SD1_SB_inst_SD1_SB_bit_inst_23_U45 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_23_n141), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_23_n140), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_23_n141), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_23_n139), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_23_n140), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_23_n138), .ZN(Feedback[47]) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_23_U44 ( .A(StateRegOutput[20]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_23_n137), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_23_n138) );
  AOI211_X1 SD1_SB_inst_SD1_SB_bit_inst_23_U43 ( .C1(
        SD1_SB_inst_SD1_SB_bit_inst_23_n136), .C2(CipherErrorVec[38]), .A(
        SD1_SB_inst_SD1_SB_bit_inst_23_n135), .B(
        SD1_SB_inst_SD1_SB_bit_inst_23_n134), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_23_n137) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_23_U42 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_23_n105), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_23_n103), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_23_n133), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_23_n134) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_23_U41 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_23_n107), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_23_n132), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_23_n131), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_23_n135) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_23_U40 ( .A1(CipherErrorVec[38]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_23_n100), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_23_n131) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_23_U39 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_23_n130), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_23_n136) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_23_U38 ( .A(StateRegOutput[22]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_23_n129), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_23_n139) );
  AOI22_X1 SD1_SB_inst_SD1_SB_bit_inst_23_U37 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_23_n128), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_23_n127), .B1(CipherErrorVec[41]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_23_n126), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_23_n129) );
  OAI211_X1 SD1_SB_inst_SD1_SB_bit_inst_23_U36 ( .C1(
        SD1_SB_inst_SD1_SB_bit_inst_23_n125), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_23_n101), .A(
        SD1_SB_inst_SD1_SB_bit_inst_23_n124), .B(
        SD1_SB_inst_SD1_SB_bit_inst_23_n123), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_23_n126) );
  NAND3_X1 SD1_SB_inst_SD1_SB_bit_inst_23_U35 ( .A1(CipherErrorVec[35]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_23_n108), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_23_n122), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_23_n123) );
  OAI22_X1 SD1_SB_inst_SD1_SB_bit_inst_23_U34 ( .A1(CipherErrorVec[38]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_23_n106), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_23_n100), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_23_n103), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_23_n122) );
  AOI22_X1 SD1_SB_inst_SD1_SB_bit_inst_23_U33 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_23_n102), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_23_n104), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_23_n105), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_23_n108), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_23_n125) );
  OAI21_X1 SD1_SB_inst_SD1_SB_bit_inst_23_U32 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_23_n100), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_23_n121), .A(
        SD1_SB_inst_SD1_SB_bit_inst_23_n120), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_23_n127) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_23_U31 ( .A(CipherErrorVec[35]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_23_n121) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_23_U30 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_23_n124), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_23_n128) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_23_U29 ( .A(StateRegOutput[21]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_23_n119), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_23_n140) );
  AOI22_X1 SD1_SB_inst_SD1_SB_bit_inst_23_U28 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_23_n105), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_23_n118), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_23_n100), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_23_n117), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_23_n119) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_23_U27 ( .A1(CipherErrorVec[38]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_23_n132), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_23_n108), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_23_n117) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_23_U26 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_23_n102), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_23_n105), .A3(CipherErrorVec[35]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_23_n132) );
  OAI22_X1 SD1_SB_inst_SD1_SB_bit_inst_23_U25 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_23_n102), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_23_n133), .B1(CipherErrorVec[41]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_23_n130), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_23_n118) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_23_U24 ( .A1(CipherErrorVec[35]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_23_n116), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_23_n133) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_23_U23 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_23_n115), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_23_n101), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_23_n116) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_23_U22 ( .A1(CipherErrorVec[38]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_23_n107), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_23_n115) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_23_U21 ( .A(StateRegOutput[23]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_23_n114), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_23_n141) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_23_U20 ( .B1(CipherErrorVec[41]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_23_n113), .A(
        SD1_SB_inst_SD1_SB_bit_inst_23_n112), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_23_n114) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_23_U19 ( .B1(CipherErrorVec[35]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_23_n124), .A(
        SD1_SB_inst_SD1_SB_bit_inst_23_n120), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_23_n112) );
  NAND3_X1 SD1_SB_inst_SD1_SB_bit_inst_23_U18 ( .A1(CipherErrorVec[38]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_23_n100), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_23_n107), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_23_n120) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_23_U17 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_23_n102), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_23_n105), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_23_n124) );
  OAI221_X1 SD1_SB_inst_SD1_SB_bit_inst_23_U16 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_23_n105), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_23_n130), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_23_n105), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_23_n111), .A(
        SD1_SB_inst_SD1_SB_bit_inst_23_n110), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_23_n113) );
  OAI21_X1 SD1_SB_inst_SD1_SB_bit_inst_23_U15 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_23_n107), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_23_n109), .A(CipherErrorVec[38]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_23_n110) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_23_U14 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_23_n102), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_23_n100), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_23_n106), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_23_n109) );
  OAI211_X1 SD1_SB_inst_SD1_SB_bit_inst_23_U13 ( .C1(CipherErrorVec[38]), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_23_n107), .A(
        SD1_SB_inst_SD1_SB_bit_inst_23_n100), .B(
        SD1_SB_inst_SD1_SB_bit_inst_23_n103), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_23_n111) );
  NAND3_X1 SD1_SB_inst_SD1_SB_bit_inst_23_U12 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_23_n102), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_23_n107), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_23_n101), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_23_n130) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_23_U11 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_23_n108), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_23_n107) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_23_U10 ( .A(CipherErrorVec[39]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_23_n106) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_23_U9 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_23_n106), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_23_n105) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_23_U8 ( .A(CipherErrorVec[38]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_23_n104) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_23_U7 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_23_n103), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_23_n102) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_23_U6 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_23_n101), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_23_n100) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_23_U5 ( .A(CipherErrorVec[37]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_23_n103) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_23_U4 ( .A(CipherErrorVec[40]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_23_n108) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_23_U3 ( .A(CipherErrorVec[36]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_23_n101) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_24_U47 ( .B1(OutputRegIn[26]), .B2(
        OutputRegIn[27]), .A(SD1_SB_inst_SD1_SB_bit_inst_24_n131), .ZN(
        Feedback[40]) );
  AOI221_X1 SD1_SB_inst_SD1_SB_bit_inst_24_U46 ( .B1(OutputRegIn[26]), .B2(
        OutputRegIn[24]), .C1(OutputRegIn[27]), .C2(OutputRegIn[24]), .A(
        OutputRegIn[25]), .ZN(SD1_SB_inst_SD1_SB_bit_inst_24_n131) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_24_U45 ( .A(StateRegOutput[27]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_24_n127), .ZN(OutputRegIn[27]) );
  AOI211_X1 SD1_SB_inst_SD1_SB_bit_inst_24_U44 ( .C1(CipherErrorVec[48]), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_24_n126), .A(
        SD1_SB_inst_SD1_SB_bit_inst_24_n125), .B(
        SD1_SB_inst_SD1_SB_bit_inst_24_n124), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_24_n127) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_24_U43 ( .A1(CipherErrorVec[42]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_24_n101), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_24_n123), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_24_n124) );
  AOI222_X1 SD1_SB_inst_SD1_SB_bit_inst_24_U42 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_24_n108), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_24_n104), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_24_n108), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_24_n122), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_24_n104), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_24_n121), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_24_n126) );
  OAI221_X1 SD1_SB_inst_SD1_SB_bit_inst_24_U41 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_24_n120), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_24_n100), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_24_n120), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_24_n102), .A(
        SD1_SB_inst_SD1_SB_bit_inst_24_n106), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_24_n121) );
  OAI211_X1 SD1_SB_inst_SD1_SB_bit_inst_24_U40 ( .C1(
        SD1_SB_inst_SD1_SB_bit_inst_24_n105), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_24_n100), .A(
        SD1_SB_inst_SD1_SB_bit_inst_24_n119), .B(
        SD1_SB_inst_SD1_SB_bit_inst_24_n102), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_24_n122) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_24_U39 ( .A(StateRegOutput[26]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_24_n118), .ZN(OutputRegIn[26]) );
  AOI211_X1 SD1_SB_inst_SD1_SB_bit_inst_24_U38 ( .C1(CipherErrorVec[48]), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_24_n117), .A(
        SD1_SB_inst_SD1_SB_bit_inst_24_n125), .B(
        SD1_SB_inst_SD1_SB_bit_inst_24_n116), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_24_n118) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_24_U37 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_24_n128), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_24_n96), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_24_n116) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_24_U36 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_24_n105), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_24_n120), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_24_n128) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_24_U35 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_24_n102), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_24_n123), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_24_n119), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_24_n125) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_24_U34 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_24_n105), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_24_n100), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_24_n119) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_24_U33 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_24_n107), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_24_n103), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_24_n123) );
  OAI22_X1 SD1_SB_inst_SD1_SB_bit_inst_24_U32 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_24_n107), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_24_n115), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_24_n114), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_24_n102), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_24_n117) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_24_U31 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_24_n100), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_24_n104), .A(
        SD1_SB_inst_SD1_SB_bit_inst_24_n105), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_24_n114) );
  AOI22_X1 SD1_SB_inst_SD1_SB_bit_inst_24_U30 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_24_n105), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_24_n100), .B1(CipherErrorVec[42]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_24_n113), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_24_n115) );
  OAI21_X1 SD1_SB_inst_SD1_SB_bit_inst_24_U29 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_24_n103), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_24_n106), .A(
        SD1_SB_inst_SD1_SB_bit_inst_24_n112), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_24_n113) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_24_U28 ( .A(StateRegOutput[24]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_24_n111), .ZN(OutputRegIn[24]) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_24_U27 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_24_n110), .B2(CipherErrorVec[44]), .A(
        SD1_SB_inst_SD1_SB_bit_inst_24_n109), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_24_n111) );
  AOI221_X1 SD1_SB_inst_SD1_SB_bit_inst_24_U26 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_24_n107), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_24_n112), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_24_n108), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_24_n129), .A(
        SD1_SB_inst_SD1_SB_bit_inst_24_n104), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_24_n109) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_24_U25 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_24_n120), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_24_n112) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_24_U24 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_24_n100), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_24_n102), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_24_n120) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_24_U23 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_24_n130), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_24_n105), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_24_n110) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_24_U22 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_24_n108), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_24_n107) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_24_U21 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_24_n106), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_24_n105) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_24_U20 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_24_n104), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_24_n103) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_24_U19 ( .A(CipherErrorVec[44]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_24_n102) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_24_U18 ( .A(CipherErrorVec[43]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_24_n101) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_24_U17 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_24_n101), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_24_n100) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_24_U16 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_24_n99), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_24_n130) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_24_U15 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_24_n97), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_24_n129) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_24_U14 ( .A(CipherErrorVec[42]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_24_n96) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_24_U13 ( .A(CipherErrorVec[47]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_24_n108) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_24_U12 ( .A(CipherErrorVec[46]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_24_n106) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_24_U11 ( .A(CipherErrorVec[45]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_24_n104) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_24_U10 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_24_n100), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_24_n107), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_24_n98) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_24_U9 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_24_n98), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_24_n104), .A(
        SD1_SB_inst_SD1_SB_bit_inst_24_n96), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_24_n99) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_24_U8 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_24_n105), .A2(CipherErrorVec[44]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_24_n95) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_24_U7 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_24_n95), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_24_n96), .A(
        SD1_SB_inst_SD1_SB_bit_inst_24_n101), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_24_n97) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_24_U6 ( .A(StateRegOutput[25]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_24_n94), .ZN(OutputRegIn[25]) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_24_U5 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_24_n107), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_24_n92), .A(
        SD1_SB_inst_SD1_SB_bit_inst_24_n93), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_24_n94) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_24_U4 ( .A1(CipherErrorVec[44]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_24_n130), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_24_n106), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_24_n93) );
  OAI22_X1 SD1_SB_inst_SD1_SB_bit_inst_24_U3 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_24_n103), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_24_n129), .B1(CipherErrorVec[48]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_24_n128), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_24_n92) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_25_U37 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_25_n110), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_25_n109), .A(
        SD1_SB_inst_SD1_SB_bit_inst_25_n108), .ZN(Feedback[41]) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_25_U36 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_25_n107), .B2(StateRegOutput[24]), .A(
        SD1_SB_inst_SD1_SB_bit_inst_25_n106), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_25_n108) );
  OAI22_X1 SD1_SB_inst_SD1_SB_bit_inst_25_U35 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_25_n109), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_25_n110), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_25_n107), .B2(StateRegOutput[24]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_25_n106) );
  AOI22_X1 SD1_SB_inst_SD1_SB_bit_inst_25_U34 ( .A1(CipherErrorVec[42]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_25_n105), .B1(CipherErrorVec[45]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_25_n104), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_25_n107) );
  OAI21_X1 SD1_SB_inst_SD1_SB_bit_inst_25_U33 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_25_n103), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_25_n102), .A(
        SD1_SB_inst_SD1_SB_bit_inst_25_n101), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_25_n104) );
  NAND3_X1 SD1_SB_inst_SD1_SB_bit_inst_25_U32 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_25_n79), .A2(CipherErrorVec[47]), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_25_n78), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_25_n101) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_25_U31 ( .A1(CipherErrorVec[42]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_25_n79), .A3(CipherErrorVec[46]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_25_n103) );
  AOI211_X1 SD1_SB_inst_SD1_SB_bit_inst_25_U30 ( .C1(
        SD1_SB_inst_SD1_SB_bit_inst_25_n100), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_25_n78), .A(CipherErrorVec[46]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_25_n80), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_25_n105) );
  XOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_25_U29 ( .A(StateRegOutput[26]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_25_n99), .Z(
        SD1_SB_inst_SD1_SB_bit_inst_25_n109) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_25_U28 ( .B1(CipherErrorVec[48]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_25_n98), .A(
        SD1_SB_inst_SD1_SB_bit_inst_25_n97), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_25_n99) );
  AOI221_X1 SD1_SB_inst_SD1_SB_bit_inst_25_U27 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_25_n77), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_25_n96), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_25_n78), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_25_n95), .A(
        SD1_SB_inst_SD1_SB_bit_inst_25_n94), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_25_n97) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_25_U26 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_25_n93), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_25_n94) );
  OAI22_X1 SD1_SB_inst_SD1_SB_bit_inst_25_U25 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_25_n92), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_25_n80), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_25_n91), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_25_n82), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_25_n98) );
  AOI211_X1 SD1_SB_inst_SD1_SB_bit_inst_25_U24 ( .C1(CipherErrorVec[42]), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_25_n100), .A(
        SD1_SB_inst_SD1_SB_bit_inst_25_n79), .B(
        SD1_SB_inst_SD1_SB_bit_inst_25_n90), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_25_n91) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_25_U23 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_25_n102), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_25_n90) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_25_U22 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_25_n77), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_25_n83), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_25_n102) );
  AOI22_X1 SD1_SB_inst_SD1_SB_bit_inst_25_U21 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_25_n77), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_25_n81), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_25_n89), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_25_n83), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_25_n92) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_25_U20 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_25_n77), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_25_n95), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_25_n89) );
  XOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_25_U19 ( .A(StateRegOutput[27]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_25_n88), .Z(
        SD1_SB_inst_SD1_SB_bit_inst_25_n110) );
  OAI21_X1 SD1_SB_inst_SD1_SB_bit_inst_25_U18 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_25_n87), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_25_n96), .A(
        SD1_SB_inst_SD1_SB_bit_inst_25_n86), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_25_n88) );
  OAI221_X1 SD1_SB_inst_SD1_SB_bit_inst_25_U17 ( .B1(CipherErrorVec[46]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_25_n85), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_25_n82), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_25_n84), .A(CipherErrorVec[48]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_25_n86) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_25_U16 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_25_n77), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_25_n79), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_25_n81), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_25_n84) );
  OAI33_X1 SD1_SB_inst_SD1_SB_bit_inst_25_U15 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_25_n79), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_25_n100), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_25_n78), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_25_n80), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_25_n83), .B3(
        SD1_SB_inst_SD1_SB_bit_inst_25_n77), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_25_n85) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_25_U14 ( .A1(CipherErrorVec[45]), .A2(
        CipherErrorVec[47]), .ZN(SD1_SB_inst_SD1_SB_bit_inst_25_n100) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_25_U13 ( .A1(CipherErrorVec[45]), .A2(
        CipherErrorVec[47]), .ZN(SD1_SB_inst_SD1_SB_bit_inst_25_n96) );
  AOI221_X1 SD1_SB_inst_SD1_SB_bit_inst_25_U12 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_25_n93), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_25_n77), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_25_n95), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_25_n77), .A(CipherErrorVec[48]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_25_n87) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_25_U11 ( .A(CipherErrorVec[42]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_25_n95) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_25_U10 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_25_n80), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_25_n82), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_25_n93) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_25_U9 ( .A(CipherErrorVec[45]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_25_n81) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_25_U8 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_25_n80), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_25_n79) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_25_U7 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_25_n78), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_25_n77) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_25_U6 ( .A(CipherErrorVec[46]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_25_n82) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_25_U5 ( .A(CipherErrorVec[47]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_25_n83) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_25_U4 ( .A(CipherErrorVec[44]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_25_n80) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_25_U3 ( .A(CipherErrorVec[43]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_25_n78) );
  OAI22_X1 SD1_SB_inst_SD1_SB_bit_inst_26_U45 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_26_n138), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_26_n137), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_26_n136), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_26_n135), .ZN(Feedback[42]) );
  XOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_26_U44 ( .A(StateRegOutput[25]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_26_n134), .Z(
        SD1_SB_inst_SD1_SB_bit_inst_26_n137) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_26_U43 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_26_n103), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_26_n133), .A(
        SD1_SB_inst_SD1_SB_bit_inst_26_n132), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_26_n134) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_26_U42 ( .A1(CipherErrorVec[45]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_26_n131), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_26_n130), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_26_n132) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_26_U41 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_26_n105), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_26_n99), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_26_n130) );
  OAI22_X1 SD1_SB_inst_SD1_SB_bit_inst_26_U40 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_26_n101), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_26_n129), .B1(CipherErrorVec[48]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_26_n128), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_26_n133) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_26_U39 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_26_n135), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_26_n136), .A(
        SD1_SB_inst_SD1_SB_bit_inst_26_n127), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_26_n138) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_26_U38 ( .A(StateRegOutput[26]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_26_n126), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_26_n127) );
  AOI211_X1 SD1_SB_inst_SD1_SB_bit_inst_26_U37 ( .C1(
        SD1_SB_inst_SD1_SB_bit_inst_26_n101), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_26_n125), .A(
        SD1_SB_inst_SD1_SB_bit_inst_26_n124), .B(
        SD1_SB_inst_SD1_SB_bit_inst_26_n123), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_26_n126) );
  AOI211_X1 SD1_SB_inst_SD1_SB_bit_inst_26_U36 ( .C1(
        SD1_SB_inst_SD1_SB_bit_inst_26_n122), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_26_n102), .A(
        SD1_SB_inst_SD1_SB_bit_inst_26_n121), .B(
        SD1_SB_inst_SD1_SB_bit_inst_26_n104), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_26_n123) );
  AOI22_X1 SD1_SB_inst_SD1_SB_bit_inst_26_U35 ( .A1(CipherErrorVec[42]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_26_n120), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_26_n99), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_26_n106), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_26_n122) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_26_U34 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_26_n102), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_26_n104), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_26_n119), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_26_n124) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_26_U33 ( .A(CipherErrorVec[48]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_26_n121) );
  OAI221_X1 SD1_SB_inst_SD1_SB_bit_inst_26_U32 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_26_n103), .B2(CipherErrorVec[48]), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_26_n103), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_26_n106), .A(CipherErrorVec[42]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_26_n118) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_26_U31 ( .A(StateRegOutput[24]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_26_n117), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_26_n136) );
  AOI22_X1 SD1_SB_inst_SD1_SB_bit_inst_26_U30 ( .A1(CipherErrorVec[45]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_26_n116), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_26_n101), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_26_n115), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_26_n117) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_26_U29 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_26_n103), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_26_n129), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_26_n115) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_26_U28 ( .A1(CipherErrorVec[42]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_26_n114), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_26_n129) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_26_U27 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_26_n120), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_26_n100), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_26_n114) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_26_U26 ( .A1(CipherErrorVec[45]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_26_n105), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_26_n120) );
  OAI21_X1 SD1_SB_inst_SD1_SB_bit_inst_26_U25 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_26_n131), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_26_n113), .A(
        SD1_SB_inst_SD1_SB_bit_inst_26_n128), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_26_n116) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_26_U24 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_26_n99), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_26_n106), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_26_n113) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_26_U23 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_26_n101), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_26_n103), .A3(CipherErrorVec[42]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_26_n131) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_26_U22 ( .A(StateRegOutput[27]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_26_n112), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_26_n135) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_26_U21 ( .B1(CipherErrorVec[48]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_26_n111), .A(
        SD1_SB_inst_SD1_SB_bit_inst_26_n110), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_26_n112) );
  AOI221_X1 SD1_SB_inst_SD1_SB_bit_inst_26_U20 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_26_n104), .B2(CipherErrorVec[42]), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_26_n102), .C2(CipherErrorVec[42]), .A(
        SD1_SB_inst_SD1_SB_bit_inst_26_n119), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_26_n110) );
  NAND3_X1 SD1_SB_inst_SD1_SB_bit_inst_26_U19 ( .A1(CipherErrorVec[45]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_26_n105), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_26_n99), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_26_n119) );
  OAI221_X1 SD1_SB_inst_SD1_SB_bit_inst_26_U18 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_26_n103), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_26_n128), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_26_n103), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_26_n109), .A(
        SD1_SB_inst_SD1_SB_bit_inst_26_n108), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_26_n111) );
  OAI21_X1 SD1_SB_inst_SD1_SB_bit_inst_26_U17 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_26_n105), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_26_n107), .A(CipherErrorVec[45]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_26_n108) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_26_U16 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_26_n101), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_26_n99), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_26_n104), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_26_n107) );
  OAI211_X1 SD1_SB_inst_SD1_SB_bit_inst_26_U15 ( .C1(CipherErrorVec[45]), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_26_n105), .A(
        SD1_SB_inst_SD1_SB_bit_inst_26_n99), .B(
        SD1_SB_inst_SD1_SB_bit_inst_26_n102), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_26_n109) );
  NAND3_X1 SD1_SB_inst_SD1_SB_bit_inst_26_U14 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_26_n101), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_26_n105), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_26_n100), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_26_n128) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_26_U13 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_26_n106), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_26_n105) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_26_U12 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_26_n104), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_26_n103) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_26_U11 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_26_n102), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_26_n101) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_26_U10 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_26_n100), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_26_n99) );
  MUX2_X1 SD1_SB_inst_SD1_SB_bit_inst_26_U9 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_26_n97), .B(
        SD1_SB_inst_SD1_SB_bit_inst_26_n98), .S(
        SD1_SB_inst_SD1_SB_bit_inst_26_n99), .Z(
        SD1_SB_inst_SD1_SB_bit_inst_26_n125) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_26_U8 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_26_n118), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_26_n97) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_26_U7 ( .A(CipherErrorVec[46]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_26_n104) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_26_U6 ( .A(CipherErrorVec[44]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_26_n102) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_26_U5 ( .A(CipherErrorVec[47]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_26_n106) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_26_U4 ( .A(CipherErrorVec[43]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_26_n100) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_26_U3 ( .A1(CipherErrorVec[45]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_26_n121), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_26_n98) );
  AOI222_X1 SD1_SB_inst_SD1_SB_bit_inst_27_U45 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_27_n141), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_27_n140), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_27_n141), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_27_n139), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_27_n140), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_27_n138), .ZN(Feedback[43]) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_27_U44 ( .A(StateRegOutput[24]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_27_n137), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_27_n138) );
  AOI211_X1 SD1_SB_inst_SD1_SB_bit_inst_27_U43 ( .C1(
        SD1_SB_inst_SD1_SB_bit_inst_27_n136), .C2(CipherErrorVec[45]), .A(
        SD1_SB_inst_SD1_SB_bit_inst_27_n135), .B(
        SD1_SB_inst_SD1_SB_bit_inst_27_n134), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_27_n137) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_27_U42 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_27_n105), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_27_n103), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_27_n133), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_27_n134) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_27_U41 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_27_n107), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_27_n132), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_27_n131), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_27_n135) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_27_U40 ( .A1(CipherErrorVec[45]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_27_n100), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_27_n131) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_27_U39 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_27_n130), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_27_n136) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_27_U38 ( .A(StateRegOutput[26]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_27_n129), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_27_n139) );
  AOI22_X1 SD1_SB_inst_SD1_SB_bit_inst_27_U37 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_27_n128), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_27_n127), .B1(CipherErrorVec[48]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_27_n126), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_27_n129) );
  OAI211_X1 SD1_SB_inst_SD1_SB_bit_inst_27_U36 ( .C1(
        SD1_SB_inst_SD1_SB_bit_inst_27_n125), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_27_n101), .A(
        SD1_SB_inst_SD1_SB_bit_inst_27_n124), .B(
        SD1_SB_inst_SD1_SB_bit_inst_27_n123), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_27_n126) );
  NAND3_X1 SD1_SB_inst_SD1_SB_bit_inst_27_U35 ( .A1(CipherErrorVec[42]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_27_n108), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_27_n122), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_27_n123) );
  OAI22_X1 SD1_SB_inst_SD1_SB_bit_inst_27_U34 ( .A1(CipherErrorVec[45]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_27_n106), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_27_n100), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_27_n103), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_27_n122) );
  AOI22_X1 SD1_SB_inst_SD1_SB_bit_inst_27_U33 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_27_n102), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_27_n104), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_27_n105), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_27_n108), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_27_n125) );
  OAI21_X1 SD1_SB_inst_SD1_SB_bit_inst_27_U32 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_27_n100), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_27_n121), .A(
        SD1_SB_inst_SD1_SB_bit_inst_27_n120), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_27_n127) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_27_U31 ( .A(CipherErrorVec[42]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_27_n121) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_27_U30 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_27_n124), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_27_n128) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_27_U29 ( .A(StateRegOutput[25]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_27_n119), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_27_n140) );
  AOI22_X1 SD1_SB_inst_SD1_SB_bit_inst_27_U28 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_27_n105), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_27_n118), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_27_n100), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_27_n117), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_27_n119) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_27_U27 ( .A1(CipherErrorVec[45]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_27_n132), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_27_n108), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_27_n117) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_27_U26 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_27_n102), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_27_n105), .A3(CipherErrorVec[42]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_27_n132) );
  OAI22_X1 SD1_SB_inst_SD1_SB_bit_inst_27_U25 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_27_n102), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_27_n133), .B1(CipherErrorVec[48]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_27_n130), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_27_n118) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_27_U24 ( .A1(CipherErrorVec[42]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_27_n116), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_27_n133) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_27_U23 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_27_n115), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_27_n101), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_27_n116) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_27_U22 ( .A1(CipherErrorVec[45]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_27_n107), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_27_n115) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_27_U21 ( .A(StateRegOutput[27]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_27_n114), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_27_n141) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_27_U20 ( .B1(CipherErrorVec[48]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_27_n113), .A(
        SD1_SB_inst_SD1_SB_bit_inst_27_n112), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_27_n114) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_27_U19 ( .B1(CipherErrorVec[42]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_27_n124), .A(
        SD1_SB_inst_SD1_SB_bit_inst_27_n120), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_27_n112) );
  NAND3_X1 SD1_SB_inst_SD1_SB_bit_inst_27_U18 ( .A1(CipherErrorVec[45]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_27_n100), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_27_n107), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_27_n120) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_27_U17 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_27_n102), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_27_n105), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_27_n124) );
  OAI221_X1 SD1_SB_inst_SD1_SB_bit_inst_27_U16 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_27_n105), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_27_n130), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_27_n105), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_27_n111), .A(
        SD1_SB_inst_SD1_SB_bit_inst_27_n110), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_27_n113) );
  OAI21_X1 SD1_SB_inst_SD1_SB_bit_inst_27_U15 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_27_n107), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_27_n109), .A(CipherErrorVec[45]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_27_n110) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_27_U14 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_27_n102), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_27_n100), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_27_n106), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_27_n109) );
  OAI211_X1 SD1_SB_inst_SD1_SB_bit_inst_27_U13 ( .C1(CipherErrorVec[45]), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_27_n107), .A(
        SD1_SB_inst_SD1_SB_bit_inst_27_n100), .B(
        SD1_SB_inst_SD1_SB_bit_inst_27_n103), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_27_n111) );
  NAND3_X1 SD1_SB_inst_SD1_SB_bit_inst_27_U12 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_27_n102), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_27_n107), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_27_n101), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_27_n130) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_27_U11 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_27_n108), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_27_n107) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_27_U10 ( .A(CipherErrorVec[46]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_27_n106) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_27_U9 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_27_n106), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_27_n105) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_27_U8 ( .A(CipherErrorVec[45]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_27_n104) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_27_U7 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_27_n103), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_27_n102) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_27_U6 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_27_n101), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_27_n100) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_27_U5 ( .A(CipherErrorVec[44]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_27_n103) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_27_U4 ( .A(CipherErrorVec[47]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_27_n108) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_27_U3 ( .A(CipherErrorVec[43]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_27_n101) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_28_U48 ( .B1(OutputRegIn[30]), .B2(
        OutputRegIn[31]), .A(SD1_SB_inst_SD1_SB_bit_inst_28_n132), .ZN(
        Feedback[36]) );
  AOI221_X1 SD1_SB_inst_SD1_SB_bit_inst_28_U47 ( .B1(OutputRegIn[30]), .B2(
        OutputRegIn[28]), .C1(OutputRegIn[31]), .C2(OutputRegIn[28]), .A(
        OutputRegIn[29]), .ZN(SD1_SB_inst_SD1_SB_bit_inst_28_n132) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_28_U46 ( .A(StateRegOutput[29]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_28_n131), .ZN(OutputRegIn[29]) );
  AOI221_X1 SD1_SB_inst_SD1_SB_bit_inst_28_U45 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_28_n130), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_28_n104), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_28_n129), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_28_n104), .A(
        SD1_SB_inst_SD1_SB_bit_inst_28_n128), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_28_n131) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_28_U44 ( .A1(CipherErrorVec[51]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_28_n103), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_28_n127), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_28_n128) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_28_U43 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_28_n100), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_28_n126), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_28_n129) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_28_U42 ( .A1(CipherErrorVec[55]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_28_n125), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_28_n130) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_28_U41 ( .A(StateRegOutput[31]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_28_n124), .ZN(OutputRegIn[31]) );
  AOI211_X1 SD1_SB_inst_SD1_SB_bit_inst_28_U40 ( .C1(CipherErrorVec[55]), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_28_n123), .A(
        SD1_SB_inst_SD1_SB_bit_inst_28_n122), .B(
        SD1_SB_inst_SD1_SB_bit_inst_28_n121), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_28_n124) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_28_U39 ( .A1(CipherErrorVec[49]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_28_n98), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_28_n120), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_28_n121) );
  AOI222_X1 SD1_SB_inst_SD1_SB_bit_inst_28_U38 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_28_n105), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_28_n101), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_28_n105), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_28_n119), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_28_n101), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_28_n118), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_28_n123) );
  OAI221_X1 SD1_SB_inst_SD1_SB_bit_inst_28_U37 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_28_n117), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_28_n97), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_28_n117), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_28_n99), .A(
        SD1_SB_inst_SD1_SB_bit_inst_28_n103), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_28_n118) );
  OAI211_X1 SD1_SB_inst_SD1_SB_bit_inst_28_U36 ( .C1(
        SD1_SB_inst_SD1_SB_bit_inst_28_n102), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_28_n97), .A(
        SD1_SB_inst_SD1_SB_bit_inst_28_n116), .B(
        SD1_SB_inst_SD1_SB_bit_inst_28_n99), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_28_n119) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_28_U35 ( .A(StateRegOutput[30]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_28_n115), .ZN(OutputRegIn[30]) );
  AOI211_X1 SD1_SB_inst_SD1_SB_bit_inst_28_U34 ( .C1(CipherErrorVec[55]), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_28_n114), .A(
        SD1_SB_inst_SD1_SB_bit_inst_28_n122), .B(
        SD1_SB_inst_SD1_SB_bit_inst_28_n113), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_28_n115) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_28_U33 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_28_n125), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_28_n93), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_28_n113) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_28_U32 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_28_n102), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_28_n117), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_28_n125) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_28_U31 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_28_n99), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_28_n120), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_28_n116), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_28_n122) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_28_U30 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_28_n102), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_28_n97), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_28_n116) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_28_U29 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_28_n104), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_28_n100), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_28_n120) );
  OAI22_X1 SD1_SB_inst_SD1_SB_bit_inst_28_U28 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_28_n104), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_28_n112), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_28_n111), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_28_n99), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_28_n114) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_28_U27 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_28_n97), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_28_n101), .A(
        SD1_SB_inst_SD1_SB_bit_inst_28_n102), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_28_n111) );
  AOI22_X1 SD1_SB_inst_SD1_SB_bit_inst_28_U26 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_28_n102), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_28_n97), .B1(CipherErrorVec[49]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_28_n110), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_28_n112) );
  OAI21_X1 SD1_SB_inst_SD1_SB_bit_inst_28_U25 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_28_n100), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_28_n103), .A(
        SD1_SB_inst_SD1_SB_bit_inst_28_n109), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_28_n110) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_28_U24 ( .A(StateRegOutput[28]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_28_n108), .ZN(OutputRegIn[28]) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_28_U23 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_28_n107), .B2(CipherErrorVec[51]), .A(
        SD1_SB_inst_SD1_SB_bit_inst_28_n106), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_28_n108) );
  AOI221_X1 SD1_SB_inst_SD1_SB_bit_inst_28_U22 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_28_n104), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_28_n109), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_28_n105), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_28_n126), .A(
        SD1_SB_inst_SD1_SB_bit_inst_28_n101), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_28_n106) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_28_U21 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_28_n117), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_28_n109) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_28_U20 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_28_n97), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_28_n99), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_28_n117) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_28_U19 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_28_n127), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_28_n102), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_28_n107) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_28_U18 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_28_n105), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_28_n104) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_28_U17 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_28_n103), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_28_n102) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_28_U16 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_28_n101), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_28_n100) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_28_U15 ( .A(CipherErrorVec[51]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_28_n99) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_28_U14 ( .A(CipherErrorVec[50]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_28_n98) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_28_U13 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_28_n98), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_28_n97) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_28_U12 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_28_n96), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_28_n127) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_28_U11 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_28_n94), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_28_n126) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_28_U10 ( .A(CipherErrorVec[49]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_28_n93) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_28_U9 ( .A(CipherErrorVec[54]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_28_n105) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_28_U8 ( .A(CipherErrorVec[53]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_28_n103) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_28_U7 ( .A(CipherErrorVec[52]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_28_n101) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_28_U6 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_28_n97), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_28_n104), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_28_n95) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_28_U5 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_28_n95), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_28_n101), .A(
        SD1_SB_inst_SD1_SB_bit_inst_28_n93), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_28_n96) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_28_U4 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_28_n102), .A2(CipherErrorVec[51]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_28_n92) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_28_U3 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_28_n92), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_28_n93), .A(
        SD1_SB_inst_SD1_SB_bit_inst_28_n98), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_28_n94) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_29_U36 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_29_n109), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_29_n108), .A(
        SD1_SB_inst_SD1_SB_bit_inst_29_n107), .ZN(Feedback[37]) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_29_U35 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_29_n106), .B2(StateRegOutput[28]), .A(
        SD1_SB_inst_SD1_SB_bit_inst_29_n105), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_29_n107) );
  OAI22_X1 SD1_SB_inst_SD1_SB_bit_inst_29_U34 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_29_n108), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_29_n109), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_29_n106), .B2(StateRegOutput[28]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_29_n105) );
  AOI22_X1 SD1_SB_inst_SD1_SB_bit_inst_29_U33 ( .A1(CipherErrorVec[49]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_29_n104), .B1(CipherErrorVec[52]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_29_n103), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_29_n106) );
  OAI21_X1 SD1_SB_inst_SD1_SB_bit_inst_29_U32 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_29_n102), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_29_n101), .A(
        SD1_SB_inst_SD1_SB_bit_inst_29_n100), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_29_n103) );
  NAND3_X1 SD1_SB_inst_SD1_SB_bit_inst_29_U31 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_29_n86), .A2(CipherErrorVec[54]), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_29_n85), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_29_n100) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_29_U30 ( .A1(CipherErrorVec[49]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_29_n86), .A3(CipherErrorVec[53]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_29_n102) );
  AOI211_X1 SD1_SB_inst_SD1_SB_bit_inst_29_U29 ( .C1(
        SD1_SB_inst_SD1_SB_bit_inst_29_n99), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_29_n85), .A(CipherErrorVec[53]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_29_n87), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_29_n104) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_29_U28 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_29_n84), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_29_n90), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_29_n101) );
  XOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_29_U27 ( .A(StateRegOutput[31]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_29_n95), .Z(
        SD1_SB_inst_SD1_SB_bit_inst_29_n109) );
  OAI21_X1 SD1_SB_inst_SD1_SB_bit_inst_29_U26 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_29_n94), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_29_n98), .A(
        SD1_SB_inst_SD1_SB_bit_inst_29_n93), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_29_n95) );
  OAI221_X1 SD1_SB_inst_SD1_SB_bit_inst_29_U25 ( .B1(CipherErrorVec[53]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_29_n92), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_29_n89), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_29_n91), .A(CipherErrorVec[55]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_29_n93) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_29_U24 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_29_n84), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_29_n86), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_29_n88), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_29_n91) );
  OAI33_X1 SD1_SB_inst_SD1_SB_bit_inst_29_U23 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_29_n86), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_29_n99), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_29_n85), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_29_n87), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_29_n90), .B3(
        SD1_SB_inst_SD1_SB_bit_inst_29_n84), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_29_n92) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_29_U22 ( .A1(CipherErrorVec[52]), .A2(
        CipherErrorVec[54]), .ZN(SD1_SB_inst_SD1_SB_bit_inst_29_n99) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_29_U21 ( .A1(CipherErrorVec[52]), .A2(
        CipherErrorVec[54]), .ZN(SD1_SB_inst_SD1_SB_bit_inst_29_n98) );
  AOI221_X1 SD1_SB_inst_SD1_SB_bit_inst_29_U20 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_29_n96), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_29_n84), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_29_n97), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_29_n84), .A(CipherErrorVec[55]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_29_n94) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_29_U19 ( .A(CipherErrorVec[49]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_29_n97) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_29_U18 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_29_n87), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_29_n89), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_29_n96) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_29_U17 ( .A(CipherErrorVec[52]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_29_n88) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_29_U16 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_29_n87), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_29_n86) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_29_U15 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_29_n85), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_29_n84) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_29_U14 ( .A(CipherErrorVec[53]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_29_n89) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_29_U13 ( .A(CipherErrorVec[54]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_29_n90) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_29_U12 ( .A(CipherErrorVec[51]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_29_n87) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_29_U11 ( .A(CipherErrorVec[50]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_29_n85) );
  XOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_29_U10 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_29_n83), .B(StateRegOutput[30]), .Z(
        SD1_SB_inst_SD1_SB_bit_inst_29_n108) );
  AOI22_X1 SD1_SB_inst_SD1_SB_bit_inst_29_U9 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_29_n77), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_29_n96), .B1(CipherErrorVec[55]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_29_n82), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_29_n83) );
  OAI22_X1 SD1_SB_inst_SD1_SB_bit_inst_29_U8 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_29_n87), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_29_n79), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_29_n89), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_29_n81), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_29_n82) );
  AOI211_X1 SD1_SB_inst_SD1_SB_bit_inst_29_U7 ( .C1(CipherErrorVec[49]), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_29_n99), .A(
        SD1_SB_inst_SD1_SB_bit_inst_29_n86), .B(
        SD1_SB_inst_SD1_SB_bit_inst_29_n80), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_29_n81) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_29_U6 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_29_n101), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_29_n80) );
  AOI22_X1 SD1_SB_inst_SD1_SB_bit_inst_29_U5 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_29_n84), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_29_n88), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_29_n90), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_29_n78), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_29_n79) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_29_U4 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_29_n84), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_29_n97), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_29_n78) );
  AOI22_X1 SD1_SB_inst_SD1_SB_bit_inst_29_U3 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_29_n84), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_29_n98), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_29_n85), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_29_n97), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_29_n77) );
  OAI22_X1 SD1_SB_inst_SD1_SB_bit_inst_30_U44 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_30_n137), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_30_n136), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_30_n135), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_30_n134), .ZN(Feedback[38]) );
  XOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_30_U43 ( .A(StateRegOutput[29]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_30_n133), .Z(
        SD1_SB_inst_SD1_SB_bit_inst_30_n136) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_30_U42 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_30_n110), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_30_n132), .A(
        SD1_SB_inst_SD1_SB_bit_inst_30_n131), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_30_n133) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_30_U41 ( .A1(CipherErrorVec[52]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_30_n130), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_30_n129), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_30_n131) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_30_U40 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_30_n112), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_30_n106), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_30_n129) );
  OAI22_X1 SD1_SB_inst_SD1_SB_bit_inst_30_U39 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_30_n108), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_30_n128), .B1(CipherErrorVec[55]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_30_n127), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_30_n132) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_30_U38 ( .A(StateRegOutput[28]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_30_n124), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_30_n135) );
  AOI22_X1 SD1_SB_inst_SD1_SB_bit_inst_30_U37 ( .A1(CipherErrorVec[52]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_30_n123), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_30_n108), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_30_n122), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_30_n124) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_30_U36 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_30_n110), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_30_n128), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_30_n122) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_30_U35 ( .A1(CipherErrorVec[49]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_30_n121), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_30_n128) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_30_U34 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_30_n126), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_30_n107), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_30_n121) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_30_U33 ( .A1(CipherErrorVec[52]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_30_n112), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_30_n126) );
  OAI21_X1 SD1_SB_inst_SD1_SB_bit_inst_30_U32 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_30_n130), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_30_n120), .A(
        SD1_SB_inst_SD1_SB_bit_inst_30_n127), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_30_n123) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_30_U31 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_30_n106), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_30_n113), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_30_n120) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_30_U30 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_30_n108), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_30_n110), .A3(CipherErrorVec[49]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_30_n130) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_30_U29 ( .A(StateRegOutput[31]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_30_n119), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_30_n134) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_30_U28 ( .B1(CipherErrorVec[55]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_30_n118), .A(
        SD1_SB_inst_SD1_SB_bit_inst_30_n117), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_30_n119) );
  AOI221_X1 SD1_SB_inst_SD1_SB_bit_inst_30_U27 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_30_n111), .B2(CipherErrorVec[49]), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_30_n109), .C2(CipherErrorVec[49]), .A(
        SD1_SB_inst_SD1_SB_bit_inst_30_n125), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_30_n117) );
  NAND3_X1 SD1_SB_inst_SD1_SB_bit_inst_30_U26 ( .A1(CipherErrorVec[52]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_30_n112), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_30_n106), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_30_n125) );
  OAI221_X1 SD1_SB_inst_SD1_SB_bit_inst_30_U25 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_30_n110), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_30_n127), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_30_n110), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_30_n116), .A(
        SD1_SB_inst_SD1_SB_bit_inst_30_n115), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_30_n118) );
  OAI21_X1 SD1_SB_inst_SD1_SB_bit_inst_30_U24 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_30_n112), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_30_n114), .A(CipherErrorVec[52]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_30_n115) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_30_U23 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_30_n108), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_30_n106), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_30_n111), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_30_n114) );
  OAI211_X1 SD1_SB_inst_SD1_SB_bit_inst_30_U22 ( .C1(CipherErrorVec[52]), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_30_n112), .A(
        SD1_SB_inst_SD1_SB_bit_inst_30_n106), .B(
        SD1_SB_inst_SD1_SB_bit_inst_30_n109), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_30_n116) );
  NAND3_X1 SD1_SB_inst_SD1_SB_bit_inst_30_U21 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_30_n108), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_30_n112), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_30_n107), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_30_n127) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_30_U20 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_30_n113), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_30_n112) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_30_U19 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_30_n111), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_30_n110) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_30_U18 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_30_n109), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_30_n108) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_30_U17 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_30_n107), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_30_n106) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_30_U16 ( .A(CipherErrorVec[53]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_30_n111) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_30_U15 ( .A(CipherErrorVec[51]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_30_n109) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_30_U14 ( .A(CipherErrorVec[54]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_30_n113) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_30_U13 ( .A(CipherErrorVec[50]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_30_n107) );
  AOI221_X1 SD1_SB_inst_SD1_SB_bit_inst_30_U12 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_30_n135), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_30_n134), .C1(StateRegOutput[30]), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_30_n104), .A(
        SD1_SB_inst_SD1_SB_bit_inst_30_n105), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_30_n137) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_30_U11 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_30_n104), .A2(StateRegOutput[30]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_30_n105) );
  AOI211_X1 SD1_SB_inst_SD1_SB_bit_inst_30_U10 ( .C1(
        SD1_SB_inst_SD1_SB_bit_inst_30_n108), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_30_n99), .A(
        SD1_SB_inst_SD1_SB_bit_inst_30_n102), .B(
        SD1_SB_inst_SD1_SB_bit_inst_30_n103), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_30_n104) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_30_U9 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_30_n111), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_30_n109), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_30_n125), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_30_n103) );
  AOI211_X1 SD1_SB_inst_SD1_SB_bit_inst_30_U8 ( .C1(
        SD1_SB_inst_SD1_SB_bit_inst_30_n109), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_30_n100), .A(
        SD1_SB_inst_SD1_SB_bit_inst_30_n111), .B(
        SD1_SB_inst_SD1_SB_bit_inst_30_n101), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_30_n102) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_30_U7 ( .A(CipherErrorVec[55]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_30_n101) );
  AOI22_X1 SD1_SB_inst_SD1_SB_bit_inst_30_U6 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_30_n106), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_30_n113), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_30_n126), .B2(CipherErrorVec[49]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_30_n100) );
  OAI22_X1 SD1_SB_inst_SD1_SB_bit_inst_30_U5 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_30_n106), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_30_n97), .B1(CipherErrorVec[52]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_30_n98), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_30_n99) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_30_U4 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_30_n106), .A2(CipherErrorVec[55]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_30_n98) );
  OAI221_X1 SD1_SB_inst_SD1_SB_bit_inst_30_U3 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_30_n110), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_30_n113), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_30_n110), .C2(CipherErrorVec[55]), .A(
        CipherErrorVec[49]), .ZN(SD1_SB_inst_SD1_SB_bit_inst_30_n97) );
  AOI222_X1 SD1_SB_inst_SD1_SB_bit_inst_31_U45 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_31_n141), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_31_n140), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_31_n141), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_31_n139), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_31_n140), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_31_n138), .ZN(Feedback[39]) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_31_U44 ( .A(StateRegOutput[28]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_31_n137), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_31_n138) );
  AOI211_X1 SD1_SB_inst_SD1_SB_bit_inst_31_U43 ( .C1(
        SD1_SB_inst_SD1_SB_bit_inst_31_n136), .C2(CipherErrorVec[52]), .A(
        SD1_SB_inst_SD1_SB_bit_inst_31_n135), .B(
        SD1_SB_inst_SD1_SB_bit_inst_31_n134), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_31_n137) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_31_U42 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_31_n105), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_31_n103), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_31_n133), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_31_n134) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_31_U41 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_31_n107), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_31_n132), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_31_n131), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_31_n135) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_31_U40 ( .A1(CipherErrorVec[52]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_31_n100), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_31_n131) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_31_U39 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_31_n130), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_31_n136) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_31_U38 ( .A(StateRegOutput[30]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_31_n129), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_31_n139) );
  AOI22_X1 SD1_SB_inst_SD1_SB_bit_inst_31_U37 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_31_n128), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_31_n127), .B1(CipherErrorVec[55]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_31_n126), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_31_n129) );
  OAI211_X1 SD1_SB_inst_SD1_SB_bit_inst_31_U36 ( .C1(
        SD1_SB_inst_SD1_SB_bit_inst_31_n125), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_31_n101), .A(
        SD1_SB_inst_SD1_SB_bit_inst_31_n124), .B(
        SD1_SB_inst_SD1_SB_bit_inst_31_n123), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_31_n126) );
  NAND3_X1 SD1_SB_inst_SD1_SB_bit_inst_31_U35 ( .A1(CipherErrorVec[49]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_31_n108), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_31_n122), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_31_n123) );
  OAI22_X1 SD1_SB_inst_SD1_SB_bit_inst_31_U34 ( .A1(CipherErrorVec[52]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_31_n106), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_31_n100), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_31_n103), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_31_n122) );
  AOI22_X1 SD1_SB_inst_SD1_SB_bit_inst_31_U33 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_31_n102), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_31_n104), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_31_n105), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_31_n108), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_31_n125) );
  OAI21_X1 SD1_SB_inst_SD1_SB_bit_inst_31_U32 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_31_n100), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_31_n121), .A(
        SD1_SB_inst_SD1_SB_bit_inst_31_n120), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_31_n127) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_31_U31 ( .A(CipherErrorVec[49]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_31_n121) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_31_U30 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_31_n124), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_31_n128) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_31_U29 ( .A(StateRegOutput[29]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_31_n119), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_31_n140) );
  AOI22_X1 SD1_SB_inst_SD1_SB_bit_inst_31_U28 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_31_n105), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_31_n118), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_31_n100), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_31_n117), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_31_n119) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_31_U27 ( .A1(CipherErrorVec[52]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_31_n132), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_31_n108), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_31_n117) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_31_U26 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_31_n102), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_31_n105), .A3(CipherErrorVec[49]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_31_n132) );
  OAI22_X1 SD1_SB_inst_SD1_SB_bit_inst_31_U25 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_31_n102), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_31_n133), .B1(CipherErrorVec[55]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_31_n130), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_31_n118) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_31_U24 ( .A1(CipherErrorVec[49]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_31_n116), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_31_n133) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_31_U23 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_31_n115), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_31_n101), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_31_n116) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_31_U22 ( .A1(CipherErrorVec[52]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_31_n107), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_31_n115) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_31_U21 ( .A(StateRegOutput[31]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_31_n114), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_31_n141) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_31_U20 ( .B1(CipherErrorVec[55]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_31_n113), .A(
        SD1_SB_inst_SD1_SB_bit_inst_31_n112), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_31_n114) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_31_U19 ( .B1(CipherErrorVec[49]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_31_n124), .A(
        SD1_SB_inst_SD1_SB_bit_inst_31_n120), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_31_n112) );
  NAND3_X1 SD1_SB_inst_SD1_SB_bit_inst_31_U18 ( .A1(CipherErrorVec[52]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_31_n100), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_31_n107), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_31_n120) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_31_U17 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_31_n102), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_31_n105), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_31_n124) );
  OAI221_X1 SD1_SB_inst_SD1_SB_bit_inst_31_U16 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_31_n105), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_31_n130), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_31_n105), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_31_n111), .A(
        SD1_SB_inst_SD1_SB_bit_inst_31_n110), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_31_n113) );
  OAI21_X1 SD1_SB_inst_SD1_SB_bit_inst_31_U15 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_31_n107), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_31_n109), .A(CipherErrorVec[52]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_31_n110) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_31_U14 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_31_n102), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_31_n100), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_31_n106), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_31_n109) );
  OAI211_X1 SD1_SB_inst_SD1_SB_bit_inst_31_U13 ( .C1(CipherErrorVec[52]), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_31_n107), .A(
        SD1_SB_inst_SD1_SB_bit_inst_31_n100), .B(
        SD1_SB_inst_SD1_SB_bit_inst_31_n103), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_31_n111) );
  NAND3_X1 SD1_SB_inst_SD1_SB_bit_inst_31_U12 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_31_n102), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_31_n107), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_31_n101), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_31_n130) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_31_U11 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_31_n108), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_31_n107) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_31_U10 ( .A(CipherErrorVec[53]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_31_n106) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_31_U9 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_31_n106), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_31_n105) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_31_U8 ( .A(CipherErrorVec[52]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_31_n104) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_31_U7 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_31_n103), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_31_n102) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_31_U6 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_31_n101), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_31_n100) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_31_U5 ( .A(CipherErrorVec[51]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_31_n103) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_31_U4 ( .A(CipherErrorVec[54]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_31_n108) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_31_U3 ( .A(CipherErrorVec[50]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_31_n101) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_32_U47 ( .B1(OutputRegIn[34]), .B2(
        OutputRegIn[35]), .A(SD1_SB_inst_SD1_SB_bit_inst_32_n131), .ZN(
        Feedback[16]) );
  AOI221_X1 SD1_SB_inst_SD1_SB_bit_inst_32_U46 ( .B1(OutputRegIn[34]), .B2(
        OutputRegIn[32]), .C1(OutputRegIn[35]), .C2(OutputRegIn[32]), .A(
        OutputRegIn[33]), .ZN(SD1_SB_inst_SD1_SB_bit_inst_32_n131) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_32_U45 ( .A(StateRegOutput[35]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_32_n127), .ZN(OutputRegIn[35]) );
  AOI211_X1 SD1_SB_inst_SD1_SB_bit_inst_32_U44 ( .C1(CipherErrorVec[62]), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_32_n126), .A(
        SD1_SB_inst_SD1_SB_bit_inst_32_n125), .B(
        SD1_SB_inst_SD1_SB_bit_inst_32_n124), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_32_n127) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_32_U43 ( .A1(CipherErrorVec[56]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_32_n101), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_32_n123), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_32_n124) );
  AOI222_X1 SD1_SB_inst_SD1_SB_bit_inst_32_U42 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_32_n108), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_32_n104), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_32_n108), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_32_n122), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_32_n104), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_32_n121), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_32_n126) );
  OAI221_X1 SD1_SB_inst_SD1_SB_bit_inst_32_U41 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_32_n120), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_32_n100), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_32_n120), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_32_n102), .A(
        SD1_SB_inst_SD1_SB_bit_inst_32_n106), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_32_n121) );
  OAI211_X1 SD1_SB_inst_SD1_SB_bit_inst_32_U40 ( .C1(
        SD1_SB_inst_SD1_SB_bit_inst_32_n105), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_32_n100), .A(
        SD1_SB_inst_SD1_SB_bit_inst_32_n119), .B(
        SD1_SB_inst_SD1_SB_bit_inst_32_n102), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_32_n122) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_32_U39 ( .A(StateRegOutput[34]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_32_n118), .ZN(OutputRegIn[34]) );
  AOI211_X1 SD1_SB_inst_SD1_SB_bit_inst_32_U38 ( .C1(CipherErrorVec[62]), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_32_n117), .A(
        SD1_SB_inst_SD1_SB_bit_inst_32_n125), .B(
        SD1_SB_inst_SD1_SB_bit_inst_32_n116), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_32_n118) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_32_U37 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_32_n128), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_32_n96), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_32_n116) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_32_U36 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_32_n105), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_32_n120), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_32_n128) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_32_U35 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_32_n102), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_32_n123), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_32_n119), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_32_n125) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_32_U34 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_32_n105), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_32_n100), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_32_n119) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_32_U33 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_32_n107), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_32_n103), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_32_n123) );
  OAI22_X1 SD1_SB_inst_SD1_SB_bit_inst_32_U32 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_32_n107), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_32_n115), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_32_n114), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_32_n102), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_32_n117) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_32_U31 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_32_n100), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_32_n104), .A(
        SD1_SB_inst_SD1_SB_bit_inst_32_n105), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_32_n114) );
  AOI22_X1 SD1_SB_inst_SD1_SB_bit_inst_32_U30 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_32_n105), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_32_n100), .B1(CipherErrorVec[56]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_32_n113), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_32_n115) );
  OAI21_X1 SD1_SB_inst_SD1_SB_bit_inst_32_U29 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_32_n103), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_32_n106), .A(
        SD1_SB_inst_SD1_SB_bit_inst_32_n112), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_32_n113) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_32_U28 ( .A(StateRegOutput[32]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_32_n111), .ZN(OutputRegIn[32]) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_32_U27 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_32_n110), .B2(CipherErrorVec[58]), .A(
        SD1_SB_inst_SD1_SB_bit_inst_32_n109), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_32_n111) );
  AOI221_X1 SD1_SB_inst_SD1_SB_bit_inst_32_U26 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_32_n107), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_32_n112), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_32_n108), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_32_n129), .A(
        SD1_SB_inst_SD1_SB_bit_inst_32_n104), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_32_n109) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_32_U25 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_32_n120), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_32_n112) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_32_U24 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_32_n100), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_32_n102), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_32_n120) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_32_U23 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_32_n130), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_32_n105), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_32_n110) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_32_U22 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_32_n108), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_32_n107) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_32_U21 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_32_n106), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_32_n105) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_32_U20 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_32_n104), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_32_n103) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_32_U19 ( .A(CipherErrorVec[58]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_32_n102) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_32_U18 ( .A(CipherErrorVec[57]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_32_n101) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_32_U17 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_32_n101), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_32_n100) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_32_U16 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_32_n99), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_32_n130) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_32_U15 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_32_n97), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_32_n129) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_32_U14 ( .A(CipherErrorVec[56]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_32_n96) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_32_U13 ( .A(CipherErrorVec[61]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_32_n108) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_32_U12 ( .A(CipherErrorVec[60]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_32_n106) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_32_U11 ( .A(CipherErrorVec[59]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_32_n104) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_32_U10 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_32_n100), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_32_n107), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_32_n98) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_32_U9 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_32_n98), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_32_n104), .A(
        SD1_SB_inst_SD1_SB_bit_inst_32_n96), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_32_n99) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_32_U8 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_32_n105), .A2(CipherErrorVec[58]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_32_n95) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_32_U7 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_32_n95), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_32_n96), .A(
        SD1_SB_inst_SD1_SB_bit_inst_32_n101), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_32_n97) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_32_U6 ( .A(StateRegOutput[33]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_32_n94), .ZN(OutputRegIn[33]) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_32_U5 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_32_n107), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_32_n92), .A(
        SD1_SB_inst_SD1_SB_bit_inst_32_n93), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_32_n94) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_32_U4 ( .A1(CipherErrorVec[58]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_32_n130), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_32_n106), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_32_n93) );
  OAI22_X1 SD1_SB_inst_SD1_SB_bit_inst_32_U3 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_32_n103), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_32_n129), .B1(CipherErrorVec[62]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_32_n128), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_32_n92) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_33_U37 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_33_n110), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_33_n109), .A(
        SD1_SB_inst_SD1_SB_bit_inst_33_n108), .ZN(Feedback[17]) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_33_U36 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_33_n107), .B2(StateRegOutput[32]), .A(
        SD1_SB_inst_SD1_SB_bit_inst_33_n106), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_33_n108) );
  OAI22_X1 SD1_SB_inst_SD1_SB_bit_inst_33_U35 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_33_n109), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_33_n110), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_33_n107), .B2(StateRegOutput[32]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_33_n106) );
  AOI22_X1 SD1_SB_inst_SD1_SB_bit_inst_33_U34 ( .A1(CipherErrorVec[56]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_33_n105), .B1(CipherErrorVec[59]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_33_n104), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_33_n107) );
  OAI21_X1 SD1_SB_inst_SD1_SB_bit_inst_33_U33 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_33_n103), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_33_n102), .A(
        SD1_SB_inst_SD1_SB_bit_inst_33_n101), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_33_n104) );
  NAND3_X1 SD1_SB_inst_SD1_SB_bit_inst_33_U32 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_33_n79), .A2(CipherErrorVec[61]), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_33_n78), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_33_n101) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_33_U31 ( .A1(CipherErrorVec[56]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_33_n79), .A3(CipherErrorVec[60]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_33_n103) );
  AOI211_X1 SD1_SB_inst_SD1_SB_bit_inst_33_U30 ( .C1(
        SD1_SB_inst_SD1_SB_bit_inst_33_n100), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_33_n78), .A(CipherErrorVec[60]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_33_n80), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_33_n105) );
  XOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_33_U29 ( .A(StateRegOutput[34]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_33_n99), .Z(
        SD1_SB_inst_SD1_SB_bit_inst_33_n109) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_33_U28 ( .B1(CipherErrorVec[62]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_33_n98), .A(
        SD1_SB_inst_SD1_SB_bit_inst_33_n97), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_33_n99) );
  AOI221_X1 SD1_SB_inst_SD1_SB_bit_inst_33_U27 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_33_n77), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_33_n96), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_33_n78), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_33_n95), .A(
        SD1_SB_inst_SD1_SB_bit_inst_33_n94), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_33_n97) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_33_U26 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_33_n93), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_33_n94) );
  OAI22_X1 SD1_SB_inst_SD1_SB_bit_inst_33_U25 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_33_n92), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_33_n80), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_33_n91), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_33_n82), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_33_n98) );
  AOI211_X1 SD1_SB_inst_SD1_SB_bit_inst_33_U24 ( .C1(CipherErrorVec[56]), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_33_n100), .A(
        SD1_SB_inst_SD1_SB_bit_inst_33_n79), .B(
        SD1_SB_inst_SD1_SB_bit_inst_33_n90), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_33_n91) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_33_U23 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_33_n102), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_33_n90) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_33_U22 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_33_n77), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_33_n83), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_33_n102) );
  AOI22_X1 SD1_SB_inst_SD1_SB_bit_inst_33_U21 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_33_n77), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_33_n81), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_33_n89), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_33_n83), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_33_n92) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_33_U20 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_33_n77), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_33_n95), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_33_n89) );
  XOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_33_U19 ( .A(StateRegOutput[35]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_33_n88), .Z(
        SD1_SB_inst_SD1_SB_bit_inst_33_n110) );
  OAI21_X1 SD1_SB_inst_SD1_SB_bit_inst_33_U18 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_33_n87), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_33_n96), .A(
        SD1_SB_inst_SD1_SB_bit_inst_33_n86), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_33_n88) );
  OAI221_X1 SD1_SB_inst_SD1_SB_bit_inst_33_U17 ( .B1(CipherErrorVec[60]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_33_n85), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_33_n82), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_33_n84), .A(CipherErrorVec[62]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_33_n86) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_33_U16 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_33_n77), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_33_n79), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_33_n81), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_33_n84) );
  OAI33_X1 SD1_SB_inst_SD1_SB_bit_inst_33_U15 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_33_n79), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_33_n100), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_33_n78), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_33_n80), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_33_n83), .B3(
        SD1_SB_inst_SD1_SB_bit_inst_33_n77), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_33_n85) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_33_U14 ( .A1(CipherErrorVec[59]), .A2(
        CipherErrorVec[61]), .ZN(SD1_SB_inst_SD1_SB_bit_inst_33_n100) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_33_U13 ( .A1(CipherErrorVec[59]), .A2(
        CipherErrorVec[61]), .ZN(SD1_SB_inst_SD1_SB_bit_inst_33_n96) );
  AOI221_X1 SD1_SB_inst_SD1_SB_bit_inst_33_U12 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_33_n93), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_33_n77), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_33_n95), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_33_n77), .A(CipherErrorVec[62]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_33_n87) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_33_U11 ( .A(CipherErrorVec[56]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_33_n95) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_33_U10 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_33_n80), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_33_n82), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_33_n93) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_33_U9 ( .A(CipherErrorVec[59]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_33_n81) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_33_U8 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_33_n80), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_33_n79) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_33_U7 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_33_n78), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_33_n77) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_33_U6 ( .A(CipherErrorVec[60]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_33_n82) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_33_U5 ( .A(CipherErrorVec[61]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_33_n83) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_33_U4 ( .A(CipherErrorVec[58]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_33_n80) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_33_U3 ( .A(CipherErrorVec[57]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_33_n78) );
  OAI22_X1 SD1_SB_inst_SD1_SB_bit_inst_34_U45 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_34_n138), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_34_n137), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_34_n136), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_34_n135), .ZN(Feedback[18]) );
  XOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_34_U44 ( .A(StateRegOutput[33]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_34_n134), .Z(
        SD1_SB_inst_SD1_SB_bit_inst_34_n137) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_34_U43 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_34_n103), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_34_n133), .A(
        SD1_SB_inst_SD1_SB_bit_inst_34_n132), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_34_n134) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_34_U42 ( .A1(CipherErrorVec[59]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_34_n131), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_34_n130), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_34_n132) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_34_U41 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_34_n105), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_34_n99), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_34_n130) );
  OAI22_X1 SD1_SB_inst_SD1_SB_bit_inst_34_U40 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_34_n101), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_34_n129), .B1(CipherErrorVec[62]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_34_n128), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_34_n133) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_34_U39 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_34_n135), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_34_n136), .A(
        SD1_SB_inst_SD1_SB_bit_inst_34_n127), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_34_n138) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_34_U38 ( .A(StateRegOutput[34]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_34_n126), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_34_n127) );
  AOI211_X1 SD1_SB_inst_SD1_SB_bit_inst_34_U37 ( .C1(
        SD1_SB_inst_SD1_SB_bit_inst_34_n101), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_34_n125), .A(
        SD1_SB_inst_SD1_SB_bit_inst_34_n124), .B(
        SD1_SB_inst_SD1_SB_bit_inst_34_n123), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_34_n126) );
  AOI211_X1 SD1_SB_inst_SD1_SB_bit_inst_34_U36 ( .C1(
        SD1_SB_inst_SD1_SB_bit_inst_34_n122), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_34_n102), .A(
        SD1_SB_inst_SD1_SB_bit_inst_34_n121), .B(
        SD1_SB_inst_SD1_SB_bit_inst_34_n104), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_34_n123) );
  AOI22_X1 SD1_SB_inst_SD1_SB_bit_inst_34_U35 ( .A1(CipherErrorVec[56]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_34_n120), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_34_n99), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_34_n106), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_34_n122) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_34_U34 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_34_n102), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_34_n104), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_34_n119), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_34_n124) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_34_U33 ( .A(CipherErrorVec[62]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_34_n121) );
  OAI221_X1 SD1_SB_inst_SD1_SB_bit_inst_34_U32 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_34_n103), .B2(CipherErrorVec[62]), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_34_n103), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_34_n106), .A(CipherErrorVec[56]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_34_n118) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_34_U31 ( .A(StateRegOutput[32]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_34_n117), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_34_n136) );
  AOI22_X1 SD1_SB_inst_SD1_SB_bit_inst_34_U30 ( .A1(CipherErrorVec[59]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_34_n116), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_34_n101), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_34_n115), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_34_n117) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_34_U29 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_34_n103), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_34_n129), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_34_n115) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_34_U28 ( .A1(CipherErrorVec[56]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_34_n114), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_34_n129) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_34_U27 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_34_n120), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_34_n100), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_34_n114) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_34_U26 ( .A1(CipherErrorVec[59]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_34_n105), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_34_n120) );
  OAI21_X1 SD1_SB_inst_SD1_SB_bit_inst_34_U25 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_34_n131), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_34_n113), .A(
        SD1_SB_inst_SD1_SB_bit_inst_34_n128), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_34_n116) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_34_U24 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_34_n99), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_34_n106), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_34_n113) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_34_U23 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_34_n101), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_34_n103), .A3(CipherErrorVec[56]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_34_n131) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_34_U22 ( .A(StateRegOutput[35]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_34_n112), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_34_n135) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_34_U21 ( .B1(CipherErrorVec[62]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_34_n111), .A(
        SD1_SB_inst_SD1_SB_bit_inst_34_n110), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_34_n112) );
  AOI221_X1 SD1_SB_inst_SD1_SB_bit_inst_34_U20 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_34_n104), .B2(CipherErrorVec[56]), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_34_n102), .C2(CipherErrorVec[56]), .A(
        SD1_SB_inst_SD1_SB_bit_inst_34_n119), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_34_n110) );
  NAND3_X1 SD1_SB_inst_SD1_SB_bit_inst_34_U19 ( .A1(CipherErrorVec[59]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_34_n105), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_34_n99), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_34_n119) );
  OAI221_X1 SD1_SB_inst_SD1_SB_bit_inst_34_U18 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_34_n103), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_34_n128), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_34_n103), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_34_n109), .A(
        SD1_SB_inst_SD1_SB_bit_inst_34_n108), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_34_n111) );
  OAI21_X1 SD1_SB_inst_SD1_SB_bit_inst_34_U17 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_34_n105), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_34_n107), .A(CipherErrorVec[59]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_34_n108) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_34_U16 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_34_n101), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_34_n99), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_34_n104), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_34_n107) );
  OAI211_X1 SD1_SB_inst_SD1_SB_bit_inst_34_U15 ( .C1(CipherErrorVec[59]), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_34_n105), .A(
        SD1_SB_inst_SD1_SB_bit_inst_34_n99), .B(
        SD1_SB_inst_SD1_SB_bit_inst_34_n102), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_34_n109) );
  NAND3_X1 SD1_SB_inst_SD1_SB_bit_inst_34_U14 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_34_n101), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_34_n105), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_34_n100), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_34_n128) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_34_U13 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_34_n106), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_34_n105) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_34_U12 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_34_n104), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_34_n103) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_34_U11 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_34_n102), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_34_n101) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_34_U10 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_34_n100), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_34_n99) );
  MUX2_X1 SD1_SB_inst_SD1_SB_bit_inst_34_U9 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_34_n97), .B(
        SD1_SB_inst_SD1_SB_bit_inst_34_n98), .S(
        SD1_SB_inst_SD1_SB_bit_inst_34_n99), .Z(
        SD1_SB_inst_SD1_SB_bit_inst_34_n125) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_34_U8 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_34_n118), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_34_n97) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_34_U7 ( .A(CipherErrorVec[60]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_34_n104) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_34_U6 ( .A(CipherErrorVec[58]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_34_n102) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_34_U5 ( .A(CipherErrorVec[61]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_34_n106) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_34_U4 ( .A(CipherErrorVec[57]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_34_n100) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_34_U3 ( .A1(CipherErrorVec[59]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_34_n121), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_34_n98) );
  AOI222_X1 SD1_SB_inst_SD1_SB_bit_inst_35_U45 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_35_n141), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_35_n140), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_35_n141), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_35_n139), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_35_n140), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_35_n138), .ZN(Feedback[19]) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_35_U44 ( .A(StateRegOutput[32]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_35_n137), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_35_n138) );
  AOI211_X1 SD1_SB_inst_SD1_SB_bit_inst_35_U43 ( .C1(
        SD1_SB_inst_SD1_SB_bit_inst_35_n136), .C2(CipherErrorVec[59]), .A(
        SD1_SB_inst_SD1_SB_bit_inst_35_n135), .B(
        SD1_SB_inst_SD1_SB_bit_inst_35_n134), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_35_n137) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_35_U42 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_35_n105), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_35_n103), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_35_n133), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_35_n134) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_35_U41 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_35_n107), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_35_n132), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_35_n131), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_35_n135) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_35_U40 ( .A1(CipherErrorVec[59]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_35_n100), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_35_n131) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_35_U39 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_35_n130), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_35_n136) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_35_U38 ( .A(StateRegOutput[34]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_35_n129), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_35_n139) );
  AOI22_X1 SD1_SB_inst_SD1_SB_bit_inst_35_U37 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_35_n128), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_35_n127), .B1(CipherErrorVec[62]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_35_n126), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_35_n129) );
  OAI211_X1 SD1_SB_inst_SD1_SB_bit_inst_35_U36 ( .C1(
        SD1_SB_inst_SD1_SB_bit_inst_35_n125), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_35_n101), .A(
        SD1_SB_inst_SD1_SB_bit_inst_35_n124), .B(
        SD1_SB_inst_SD1_SB_bit_inst_35_n123), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_35_n126) );
  NAND3_X1 SD1_SB_inst_SD1_SB_bit_inst_35_U35 ( .A1(CipherErrorVec[56]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_35_n108), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_35_n122), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_35_n123) );
  OAI22_X1 SD1_SB_inst_SD1_SB_bit_inst_35_U34 ( .A1(CipherErrorVec[59]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_35_n106), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_35_n100), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_35_n103), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_35_n122) );
  AOI22_X1 SD1_SB_inst_SD1_SB_bit_inst_35_U33 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_35_n102), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_35_n104), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_35_n105), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_35_n108), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_35_n125) );
  OAI21_X1 SD1_SB_inst_SD1_SB_bit_inst_35_U32 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_35_n100), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_35_n121), .A(
        SD1_SB_inst_SD1_SB_bit_inst_35_n120), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_35_n127) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_35_U31 ( .A(CipherErrorVec[56]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_35_n121) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_35_U30 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_35_n124), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_35_n128) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_35_U29 ( .A(StateRegOutput[33]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_35_n119), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_35_n140) );
  AOI22_X1 SD1_SB_inst_SD1_SB_bit_inst_35_U28 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_35_n105), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_35_n118), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_35_n100), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_35_n117), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_35_n119) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_35_U27 ( .A1(CipherErrorVec[59]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_35_n132), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_35_n108), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_35_n117) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_35_U26 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_35_n102), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_35_n105), .A3(CipherErrorVec[56]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_35_n132) );
  OAI22_X1 SD1_SB_inst_SD1_SB_bit_inst_35_U25 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_35_n102), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_35_n133), .B1(CipherErrorVec[62]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_35_n130), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_35_n118) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_35_U24 ( .A1(CipherErrorVec[56]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_35_n116), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_35_n133) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_35_U23 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_35_n115), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_35_n101), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_35_n116) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_35_U22 ( .A1(CipherErrorVec[59]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_35_n107), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_35_n115) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_35_U21 ( .A(StateRegOutput[35]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_35_n114), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_35_n141) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_35_U20 ( .B1(CipherErrorVec[62]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_35_n113), .A(
        SD1_SB_inst_SD1_SB_bit_inst_35_n112), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_35_n114) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_35_U19 ( .B1(CipherErrorVec[56]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_35_n124), .A(
        SD1_SB_inst_SD1_SB_bit_inst_35_n120), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_35_n112) );
  NAND3_X1 SD1_SB_inst_SD1_SB_bit_inst_35_U18 ( .A1(CipherErrorVec[59]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_35_n100), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_35_n107), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_35_n120) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_35_U17 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_35_n102), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_35_n105), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_35_n124) );
  OAI221_X1 SD1_SB_inst_SD1_SB_bit_inst_35_U16 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_35_n105), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_35_n130), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_35_n105), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_35_n111), .A(
        SD1_SB_inst_SD1_SB_bit_inst_35_n110), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_35_n113) );
  OAI21_X1 SD1_SB_inst_SD1_SB_bit_inst_35_U15 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_35_n107), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_35_n109), .A(CipherErrorVec[59]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_35_n110) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_35_U14 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_35_n102), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_35_n100), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_35_n106), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_35_n109) );
  OAI211_X1 SD1_SB_inst_SD1_SB_bit_inst_35_U13 ( .C1(CipherErrorVec[59]), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_35_n107), .A(
        SD1_SB_inst_SD1_SB_bit_inst_35_n100), .B(
        SD1_SB_inst_SD1_SB_bit_inst_35_n103), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_35_n111) );
  NAND3_X1 SD1_SB_inst_SD1_SB_bit_inst_35_U12 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_35_n102), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_35_n107), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_35_n101), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_35_n130) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_35_U11 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_35_n108), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_35_n107) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_35_U10 ( .A(CipherErrorVec[60]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_35_n106) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_35_U9 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_35_n106), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_35_n105) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_35_U8 ( .A(CipherErrorVec[59]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_35_n104) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_35_U7 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_35_n103), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_35_n102) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_35_U6 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_35_n101), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_35_n100) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_35_U5 ( .A(CipherErrorVec[58]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_35_n103) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_35_U4 ( .A(CipherErrorVec[61]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_35_n108) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_35_U3 ( .A(CipherErrorVec[57]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_35_n101) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_36_U47 ( .B1(OutputRegIn[38]), .B2(
        OutputRegIn[39]), .A(SD1_SB_inst_SD1_SB_bit_inst_36_n131), .ZN(
        Feedback[28]) );
  AOI221_X1 SD1_SB_inst_SD1_SB_bit_inst_36_U46 ( .B1(OutputRegIn[38]), .B2(
        OutputRegIn[36]), .C1(OutputRegIn[39]), .C2(OutputRegIn[36]), .A(
        OutputRegIn[37]), .ZN(SD1_SB_inst_SD1_SB_bit_inst_36_n131) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_36_U45 ( .A(StateRegOutput[39]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_36_n127), .ZN(OutputRegIn[39]) );
  AOI211_X1 SD1_SB_inst_SD1_SB_bit_inst_36_U44 ( .C1(CipherErrorVec[69]), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_36_n126), .A(
        SD1_SB_inst_SD1_SB_bit_inst_36_n125), .B(
        SD1_SB_inst_SD1_SB_bit_inst_36_n124), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_36_n127) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_36_U43 ( .A1(CipherErrorVec[63]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_36_n101), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_36_n123), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_36_n124) );
  AOI222_X1 SD1_SB_inst_SD1_SB_bit_inst_36_U42 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_36_n108), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_36_n104), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_36_n108), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_36_n122), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_36_n104), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_36_n121), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_36_n126) );
  OAI221_X1 SD1_SB_inst_SD1_SB_bit_inst_36_U41 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_36_n120), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_36_n100), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_36_n120), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_36_n102), .A(
        SD1_SB_inst_SD1_SB_bit_inst_36_n106), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_36_n121) );
  OAI211_X1 SD1_SB_inst_SD1_SB_bit_inst_36_U40 ( .C1(
        SD1_SB_inst_SD1_SB_bit_inst_36_n105), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_36_n100), .A(
        SD1_SB_inst_SD1_SB_bit_inst_36_n119), .B(
        SD1_SB_inst_SD1_SB_bit_inst_36_n102), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_36_n122) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_36_U39 ( .A(StateRegOutput[38]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_36_n118), .ZN(OutputRegIn[38]) );
  AOI211_X1 SD1_SB_inst_SD1_SB_bit_inst_36_U38 ( .C1(CipherErrorVec[69]), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_36_n117), .A(
        SD1_SB_inst_SD1_SB_bit_inst_36_n125), .B(
        SD1_SB_inst_SD1_SB_bit_inst_36_n116), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_36_n118) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_36_U37 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_36_n128), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_36_n96), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_36_n116) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_36_U36 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_36_n105), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_36_n120), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_36_n128) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_36_U35 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_36_n102), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_36_n123), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_36_n119), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_36_n125) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_36_U34 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_36_n105), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_36_n100), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_36_n119) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_36_U33 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_36_n107), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_36_n103), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_36_n123) );
  OAI22_X1 SD1_SB_inst_SD1_SB_bit_inst_36_U32 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_36_n107), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_36_n115), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_36_n114), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_36_n102), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_36_n117) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_36_U31 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_36_n100), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_36_n104), .A(
        SD1_SB_inst_SD1_SB_bit_inst_36_n105), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_36_n114) );
  AOI22_X1 SD1_SB_inst_SD1_SB_bit_inst_36_U30 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_36_n105), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_36_n100), .B1(CipherErrorVec[63]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_36_n113), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_36_n115) );
  OAI21_X1 SD1_SB_inst_SD1_SB_bit_inst_36_U29 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_36_n103), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_36_n106), .A(
        SD1_SB_inst_SD1_SB_bit_inst_36_n112), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_36_n113) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_36_U28 ( .A(StateRegOutput[36]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_36_n111), .ZN(OutputRegIn[36]) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_36_U27 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_36_n110), .B2(CipherErrorVec[65]), .A(
        SD1_SB_inst_SD1_SB_bit_inst_36_n109), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_36_n111) );
  AOI221_X1 SD1_SB_inst_SD1_SB_bit_inst_36_U26 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_36_n107), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_36_n112), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_36_n108), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_36_n129), .A(
        SD1_SB_inst_SD1_SB_bit_inst_36_n104), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_36_n109) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_36_U25 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_36_n120), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_36_n112) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_36_U24 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_36_n100), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_36_n102), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_36_n120) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_36_U23 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_36_n130), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_36_n105), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_36_n110) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_36_U22 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_36_n108), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_36_n107) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_36_U21 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_36_n106), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_36_n105) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_36_U20 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_36_n104), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_36_n103) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_36_U19 ( .A(CipherErrorVec[65]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_36_n102) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_36_U18 ( .A(CipherErrorVec[64]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_36_n101) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_36_U17 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_36_n101), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_36_n100) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_36_U16 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_36_n99), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_36_n130) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_36_U15 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_36_n97), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_36_n129) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_36_U14 ( .A(CipherErrorVec[63]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_36_n96) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_36_U13 ( .A(CipherErrorVec[68]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_36_n108) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_36_U12 ( .A(CipherErrorVec[67]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_36_n106) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_36_U11 ( .A(CipherErrorVec[66]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_36_n104) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_36_U10 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_36_n100), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_36_n107), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_36_n98) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_36_U9 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_36_n98), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_36_n104), .A(
        SD1_SB_inst_SD1_SB_bit_inst_36_n96), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_36_n99) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_36_U8 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_36_n105), .A2(CipherErrorVec[65]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_36_n95) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_36_U7 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_36_n95), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_36_n96), .A(
        SD1_SB_inst_SD1_SB_bit_inst_36_n101), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_36_n97) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_36_U6 ( .A(StateRegOutput[37]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_36_n94), .ZN(OutputRegIn[37]) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_36_U5 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_36_n107), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_36_n92), .A(
        SD1_SB_inst_SD1_SB_bit_inst_36_n93), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_36_n94) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_36_U4 ( .A1(CipherErrorVec[65]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_36_n130), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_36_n106), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_36_n93) );
  OAI22_X1 SD1_SB_inst_SD1_SB_bit_inst_36_U3 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_36_n103), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_36_n129), .B1(CipherErrorVec[69]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_36_n128), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_36_n92) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_37_U37 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_37_n110), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_37_n109), .A(
        SD1_SB_inst_SD1_SB_bit_inst_37_n108), .ZN(Feedback[29]) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_37_U36 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_37_n107), .B2(StateRegOutput[36]), .A(
        SD1_SB_inst_SD1_SB_bit_inst_37_n106), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_37_n108) );
  OAI22_X1 SD1_SB_inst_SD1_SB_bit_inst_37_U35 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_37_n109), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_37_n110), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_37_n107), .B2(StateRegOutput[36]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_37_n106) );
  AOI22_X1 SD1_SB_inst_SD1_SB_bit_inst_37_U34 ( .A1(CipherErrorVec[63]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_37_n105), .B1(CipherErrorVec[66]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_37_n104), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_37_n107) );
  OAI21_X1 SD1_SB_inst_SD1_SB_bit_inst_37_U33 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_37_n103), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_37_n102), .A(
        SD1_SB_inst_SD1_SB_bit_inst_37_n101), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_37_n104) );
  NAND3_X1 SD1_SB_inst_SD1_SB_bit_inst_37_U32 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_37_n79), .A2(CipherErrorVec[68]), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_37_n78), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_37_n101) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_37_U31 ( .A1(CipherErrorVec[63]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_37_n79), .A3(CipherErrorVec[67]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_37_n103) );
  AOI211_X1 SD1_SB_inst_SD1_SB_bit_inst_37_U30 ( .C1(
        SD1_SB_inst_SD1_SB_bit_inst_37_n100), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_37_n78), .A(CipherErrorVec[67]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_37_n80), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_37_n105) );
  XOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_37_U29 ( .A(StateRegOutput[38]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_37_n99), .Z(
        SD1_SB_inst_SD1_SB_bit_inst_37_n109) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_37_U28 ( .B1(CipherErrorVec[69]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_37_n98), .A(
        SD1_SB_inst_SD1_SB_bit_inst_37_n97), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_37_n99) );
  AOI221_X1 SD1_SB_inst_SD1_SB_bit_inst_37_U27 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_37_n77), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_37_n96), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_37_n78), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_37_n95), .A(
        SD1_SB_inst_SD1_SB_bit_inst_37_n94), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_37_n97) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_37_U26 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_37_n93), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_37_n94) );
  OAI22_X1 SD1_SB_inst_SD1_SB_bit_inst_37_U25 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_37_n92), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_37_n80), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_37_n91), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_37_n82), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_37_n98) );
  AOI211_X1 SD1_SB_inst_SD1_SB_bit_inst_37_U24 ( .C1(CipherErrorVec[63]), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_37_n100), .A(
        SD1_SB_inst_SD1_SB_bit_inst_37_n79), .B(
        SD1_SB_inst_SD1_SB_bit_inst_37_n90), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_37_n91) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_37_U23 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_37_n102), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_37_n90) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_37_U22 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_37_n77), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_37_n83), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_37_n102) );
  AOI22_X1 SD1_SB_inst_SD1_SB_bit_inst_37_U21 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_37_n77), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_37_n81), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_37_n89), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_37_n83), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_37_n92) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_37_U20 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_37_n77), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_37_n95), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_37_n89) );
  XOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_37_U19 ( .A(StateRegOutput[39]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_37_n88), .Z(
        SD1_SB_inst_SD1_SB_bit_inst_37_n110) );
  OAI21_X1 SD1_SB_inst_SD1_SB_bit_inst_37_U18 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_37_n87), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_37_n96), .A(
        SD1_SB_inst_SD1_SB_bit_inst_37_n86), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_37_n88) );
  OAI221_X1 SD1_SB_inst_SD1_SB_bit_inst_37_U17 ( .B1(CipherErrorVec[67]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_37_n85), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_37_n82), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_37_n84), .A(CipherErrorVec[69]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_37_n86) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_37_U16 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_37_n77), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_37_n79), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_37_n81), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_37_n84) );
  OAI33_X1 SD1_SB_inst_SD1_SB_bit_inst_37_U15 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_37_n79), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_37_n100), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_37_n78), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_37_n80), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_37_n83), .B3(
        SD1_SB_inst_SD1_SB_bit_inst_37_n77), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_37_n85) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_37_U14 ( .A1(CipherErrorVec[66]), .A2(
        CipherErrorVec[68]), .ZN(SD1_SB_inst_SD1_SB_bit_inst_37_n100) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_37_U13 ( .A1(CipherErrorVec[66]), .A2(
        CipherErrorVec[68]), .ZN(SD1_SB_inst_SD1_SB_bit_inst_37_n96) );
  AOI221_X1 SD1_SB_inst_SD1_SB_bit_inst_37_U12 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_37_n93), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_37_n77), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_37_n95), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_37_n77), .A(CipherErrorVec[69]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_37_n87) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_37_U11 ( .A(CipherErrorVec[63]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_37_n95) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_37_U10 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_37_n80), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_37_n82), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_37_n93) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_37_U9 ( .A(CipherErrorVec[66]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_37_n81) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_37_U8 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_37_n80), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_37_n79) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_37_U7 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_37_n78), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_37_n77) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_37_U6 ( .A(CipherErrorVec[67]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_37_n82) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_37_U5 ( .A(CipherErrorVec[68]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_37_n83) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_37_U4 ( .A(CipherErrorVec[65]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_37_n80) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_37_U3 ( .A(CipherErrorVec[64]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_37_n78) );
  OAI22_X1 SD1_SB_inst_SD1_SB_bit_inst_38_U45 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_38_n138), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_38_n137), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_38_n136), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_38_n135), .ZN(Feedback[30]) );
  XOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_38_U44 ( .A(StateRegOutput[37]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_38_n134), .Z(
        SD1_SB_inst_SD1_SB_bit_inst_38_n137) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_38_U43 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_38_n103), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_38_n133), .A(
        SD1_SB_inst_SD1_SB_bit_inst_38_n132), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_38_n134) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_38_U42 ( .A1(CipherErrorVec[66]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_38_n131), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_38_n130), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_38_n132) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_38_U41 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_38_n105), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_38_n99), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_38_n130) );
  OAI22_X1 SD1_SB_inst_SD1_SB_bit_inst_38_U40 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_38_n101), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_38_n129), .B1(CipherErrorVec[69]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_38_n128), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_38_n133) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_38_U39 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_38_n135), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_38_n136), .A(
        SD1_SB_inst_SD1_SB_bit_inst_38_n127), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_38_n138) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_38_U38 ( .A(StateRegOutput[38]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_38_n126), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_38_n127) );
  AOI211_X1 SD1_SB_inst_SD1_SB_bit_inst_38_U37 ( .C1(
        SD1_SB_inst_SD1_SB_bit_inst_38_n101), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_38_n125), .A(
        SD1_SB_inst_SD1_SB_bit_inst_38_n124), .B(
        SD1_SB_inst_SD1_SB_bit_inst_38_n123), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_38_n126) );
  AOI211_X1 SD1_SB_inst_SD1_SB_bit_inst_38_U36 ( .C1(
        SD1_SB_inst_SD1_SB_bit_inst_38_n122), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_38_n102), .A(
        SD1_SB_inst_SD1_SB_bit_inst_38_n121), .B(
        SD1_SB_inst_SD1_SB_bit_inst_38_n104), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_38_n123) );
  AOI22_X1 SD1_SB_inst_SD1_SB_bit_inst_38_U35 ( .A1(CipherErrorVec[63]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_38_n120), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_38_n99), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_38_n106), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_38_n122) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_38_U34 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_38_n102), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_38_n104), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_38_n119), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_38_n124) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_38_U33 ( .A(CipherErrorVec[69]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_38_n121) );
  OAI221_X1 SD1_SB_inst_SD1_SB_bit_inst_38_U32 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_38_n103), .B2(CipherErrorVec[69]), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_38_n103), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_38_n106), .A(CipherErrorVec[63]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_38_n118) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_38_U31 ( .A(StateRegOutput[36]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_38_n117), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_38_n136) );
  AOI22_X1 SD1_SB_inst_SD1_SB_bit_inst_38_U30 ( .A1(CipherErrorVec[66]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_38_n116), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_38_n101), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_38_n115), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_38_n117) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_38_U29 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_38_n103), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_38_n129), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_38_n115) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_38_U28 ( .A1(CipherErrorVec[63]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_38_n114), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_38_n129) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_38_U27 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_38_n120), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_38_n100), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_38_n114) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_38_U26 ( .A1(CipherErrorVec[66]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_38_n105), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_38_n120) );
  OAI21_X1 SD1_SB_inst_SD1_SB_bit_inst_38_U25 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_38_n131), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_38_n113), .A(
        SD1_SB_inst_SD1_SB_bit_inst_38_n128), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_38_n116) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_38_U24 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_38_n99), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_38_n106), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_38_n113) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_38_U23 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_38_n101), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_38_n103), .A3(CipherErrorVec[63]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_38_n131) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_38_U22 ( .A(StateRegOutput[39]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_38_n112), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_38_n135) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_38_U21 ( .B1(CipherErrorVec[69]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_38_n111), .A(
        SD1_SB_inst_SD1_SB_bit_inst_38_n110), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_38_n112) );
  AOI221_X1 SD1_SB_inst_SD1_SB_bit_inst_38_U20 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_38_n104), .B2(CipherErrorVec[63]), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_38_n102), .C2(CipherErrorVec[63]), .A(
        SD1_SB_inst_SD1_SB_bit_inst_38_n119), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_38_n110) );
  NAND3_X1 SD1_SB_inst_SD1_SB_bit_inst_38_U19 ( .A1(CipherErrorVec[66]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_38_n105), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_38_n99), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_38_n119) );
  OAI221_X1 SD1_SB_inst_SD1_SB_bit_inst_38_U18 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_38_n103), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_38_n128), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_38_n103), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_38_n109), .A(
        SD1_SB_inst_SD1_SB_bit_inst_38_n108), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_38_n111) );
  OAI21_X1 SD1_SB_inst_SD1_SB_bit_inst_38_U17 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_38_n105), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_38_n107), .A(CipherErrorVec[66]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_38_n108) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_38_U16 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_38_n101), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_38_n99), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_38_n104), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_38_n107) );
  OAI211_X1 SD1_SB_inst_SD1_SB_bit_inst_38_U15 ( .C1(CipherErrorVec[66]), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_38_n105), .A(
        SD1_SB_inst_SD1_SB_bit_inst_38_n99), .B(
        SD1_SB_inst_SD1_SB_bit_inst_38_n102), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_38_n109) );
  NAND3_X1 SD1_SB_inst_SD1_SB_bit_inst_38_U14 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_38_n101), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_38_n105), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_38_n100), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_38_n128) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_38_U13 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_38_n106), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_38_n105) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_38_U12 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_38_n104), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_38_n103) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_38_U11 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_38_n102), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_38_n101) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_38_U10 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_38_n100), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_38_n99) );
  MUX2_X1 SD1_SB_inst_SD1_SB_bit_inst_38_U9 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_38_n97), .B(
        SD1_SB_inst_SD1_SB_bit_inst_38_n98), .S(
        SD1_SB_inst_SD1_SB_bit_inst_38_n99), .Z(
        SD1_SB_inst_SD1_SB_bit_inst_38_n125) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_38_U8 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_38_n118), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_38_n97) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_38_U7 ( .A(CipherErrorVec[67]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_38_n104) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_38_U6 ( .A(CipherErrorVec[65]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_38_n102) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_38_U5 ( .A(CipherErrorVec[68]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_38_n106) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_38_U4 ( .A(CipherErrorVec[64]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_38_n100) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_38_U3 ( .A1(CipherErrorVec[66]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_38_n121), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_38_n98) );
  AOI222_X1 SD1_SB_inst_SD1_SB_bit_inst_39_U45 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_39_n141), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_39_n140), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_39_n141), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_39_n139), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_39_n140), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_39_n138), .ZN(Feedback[31]) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_39_U44 ( .A(StateRegOutput[36]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_39_n137), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_39_n138) );
  AOI211_X1 SD1_SB_inst_SD1_SB_bit_inst_39_U43 ( .C1(
        SD1_SB_inst_SD1_SB_bit_inst_39_n136), .C2(CipherErrorVec[66]), .A(
        SD1_SB_inst_SD1_SB_bit_inst_39_n135), .B(
        SD1_SB_inst_SD1_SB_bit_inst_39_n134), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_39_n137) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_39_U42 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_39_n105), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_39_n103), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_39_n133), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_39_n134) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_39_U41 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_39_n107), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_39_n132), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_39_n131), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_39_n135) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_39_U40 ( .A1(CipherErrorVec[66]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_39_n100), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_39_n131) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_39_U39 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_39_n130), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_39_n136) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_39_U38 ( .A(StateRegOutput[38]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_39_n129), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_39_n139) );
  AOI22_X1 SD1_SB_inst_SD1_SB_bit_inst_39_U37 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_39_n128), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_39_n127), .B1(CipherErrorVec[69]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_39_n126), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_39_n129) );
  OAI211_X1 SD1_SB_inst_SD1_SB_bit_inst_39_U36 ( .C1(
        SD1_SB_inst_SD1_SB_bit_inst_39_n125), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_39_n101), .A(
        SD1_SB_inst_SD1_SB_bit_inst_39_n124), .B(
        SD1_SB_inst_SD1_SB_bit_inst_39_n123), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_39_n126) );
  NAND3_X1 SD1_SB_inst_SD1_SB_bit_inst_39_U35 ( .A1(CipherErrorVec[63]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_39_n108), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_39_n122), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_39_n123) );
  OAI22_X1 SD1_SB_inst_SD1_SB_bit_inst_39_U34 ( .A1(CipherErrorVec[66]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_39_n106), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_39_n100), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_39_n103), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_39_n122) );
  AOI22_X1 SD1_SB_inst_SD1_SB_bit_inst_39_U33 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_39_n102), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_39_n104), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_39_n105), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_39_n108), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_39_n125) );
  OAI21_X1 SD1_SB_inst_SD1_SB_bit_inst_39_U32 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_39_n100), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_39_n121), .A(
        SD1_SB_inst_SD1_SB_bit_inst_39_n120), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_39_n127) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_39_U31 ( .A(CipherErrorVec[63]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_39_n121) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_39_U30 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_39_n124), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_39_n128) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_39_U29 ( .A(StateRegOutput[37]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_39_n119), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_39_n140) );
  AOI22_X1 SD1_SB_inst_SD1_SB_bit_inst_39_U28 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_39_n105), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_39_n118), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_39_n100), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_39_n117), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_39_n119) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_39_U27 ( .A1(CipherErrorVec[66]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_39_n132), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_39_n108), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_39_n117) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_39_U26 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_39_n102), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_39_n105), .A3(CipherErrorVec[63]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_39_n132) );
  OAI22_X1 SD1_SB_inst_SD1_SB_bit_inst_39_U25 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_39_n102), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_39_n133), .B1(CipherErrorVec[69]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_39_n130), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_39_n118) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_39_U24 ( .A1(CipherErrorVec[63]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_39_n116), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_39_n133) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_39_U23 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_39_n115), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_39_n101), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_39_n116) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_39_U22 ( .A1(CipherErrorVec[66]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_39_n107), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_39_n115) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_39_U21 ( .A(StateRegOutput[39]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_39_n114), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_39_n141) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_39_U20 ( .B1(CipherErrorVec[69]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_39_n113), .A(
        SD1_SB_inst_SD1_SB_bit_inst_39_n112), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_39_n114) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_39_U19 ( .B1(CipherErrorVec[63]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_39_n124), .A(
        SD1_SB_inst_SD1_SB_bit_inst_39_n120), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_39_n112) );
  NAND3_X1 SD1_SB_inst_SD1_SB_bit_inst_39_U18 ( .A1(CipherErrorVec[66]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_39_n100), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_39_n107), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_39_n120) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_39_U17 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_39_n102), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_39_n105), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_39_n124) );
  OAI221_X1 SD1_SB_inst_SD1_SB_bit_inst_39_U16 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_39_n105), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_39_n130), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_39_n105), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_39_n111), .A(
        SD1_SB_inst_SD1_SB_bit_inst_39_n110), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_39_n113) );
  OAI21_X1 SD1_SB_inst_SD1_SB_bit_inst_39_U15 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_39_n107), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_39_n109), .A(CipherErrorVec[66]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_39_n110) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_39_U14 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_39_n102), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_39_n100), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_39_n106), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_39_n109) );
  OAI211_X1 SD1_SB_inst_SD1_SB_bit_inst_39_U13 ( .C1(CipherErrorVec[66]), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_39_n107), .A(
        SD1_SB_inst_SD1_SB_bit_inst_39_n100), .B(
        SD1_SB_inst_SD1_SB_bit_inst_39_n103), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_39_n111) );
  NAND3_X1 SD1_SB_inst_SD1_SB_bit_inst_39_U12 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_39_n102), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_39_n107), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_39_n101), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_39_n130) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_39_U11 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_39_n108), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_39_n107) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_39_U10 ( .A(CipherErrorVec[67]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_39_n106) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_39_U9 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_39_n106), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_39_n105) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_39_U8 ( .A(CipherErrorVec[66]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_39_n104) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_39_U7 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_39_n103), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_39_n102) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_39_U6 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_39_n101), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_39_n100) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_39_U5 ( .A(CipherErrorVec[65]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_39_n103) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_39_U4 ( .A(CipherErrorVec[68]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_39_n108) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_39_U3 ( .A(CipherErrorVec[64]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_39_n101) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_40_U47 ( .B1(OutputRegIn[42]), .B2(
        OutputRegIn[43]), .A(SD1_SB_inst_SD1_SB_bit_inst_40_n131), .ZN(
        Feedback[24]) );
  AOI221_X1 SD1_SB_inst_SD1_SB_bit_inst_40_U46 ( .B1(OutputRegIn[42]), .B2(
        OutputRegIn[40]), .C1(OutputRegIn[43]), .C2(OutputRegIn[40]), .A(
        OutputRegIn[41]), .ZN(SD1_SB_inst_SD1_SB_bit_inst_40_n131) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_40_U45 ( .A(StateRegOutput[43]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_40_n127), .ZN(OutputRegIn[43]) );
  AOI211_X1 SD1_SB_inst_SD1_SB_bit_inst_40_U44 ( .C1(CipherErrorVec[76]), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_40_n126), .A(
        SD1_SB_inst_SD1_SB_bit_inst_40_n125), .B(
        SD1_SB_inst_SD1_SB_bit_inst_40_n124), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_40_n127) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_40_U43 ( .A1(CipherErrorVec[70]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_40_n101), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_40_n123), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_40_n124) );
  AOI222_X1 SD1_SB_inst_SD1_SB_bit_inst_40_U42 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_40_n108), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_40_n104), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_40_n108), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_40_n122), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_40_n104), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_40_n121), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_40_n126) );
  OAI221_X1 SD1_SB_inst_SD1_SB_bit_inst_40_U41 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_40_n120), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_40_n100), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_40_n120), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_40_n102), .A(
        SD1_SB_inst_SD1_SB_bit_inst_40_n106), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_40_n121) );
  OAI211_X1 SD1_SB_inst_SD1_SB_bit_inst_40_U40 ( .C1(
        SD1_SB_inst_SD1_SB_bit_inst_40_n105), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_40_n100), .A(
        SD1_SB_inst_SD1_SB_bit_inst_40_n119), .B(
        SD1_SB_inst_SD1_SB_bit_inst_40_n102), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_40_n122) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_40_U39 ( .A(StateRegOutput[42]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_40_n118), .ZN(OutputRegIn[42]) );
  AOI211_X1 SD1_SB_inst_SD1_SB_bit_inst_40_U38 ( .C1(CipherErrorVec[76]), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_40_n117), .A(
        SD1_SB_inst_SD1_SB_bit_inst_40_n125), .B(
        SD1_SB_inst_SD1_SB_bit_inst_40_n116), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_40_n118) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_40_U37 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_40_n128), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_40_n96), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_40_n116) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_40_U36 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_40_n105), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_40_n120), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_40_n128) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_40_U35 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_40_n102), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_40_n123), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_40_n119), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_40_n125) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_40_U34 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_40_n105), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_40_n100), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_40_n119) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_40_U33 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_40_n107), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_40_n103), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_40_n123) );
  OAI22_X1 SD1_SB_inst_SD1_SB_bit_inst_40_U32 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_40_n107), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_40_n115), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_40_n114), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_40_n102), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_40_n117) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_40_U31 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_40_n100), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_40_n104), .A(
        SD1_SB_inst_SD1_SB_bit_inst_40_n105), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_40_n114) );
  AOI22_X1 SD1_SB_inst_SD1_SB_bit_inst_40_U30 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_40_n105), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_40_n100), .B1(CipherErrorVec[70]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_40_n113), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_40_n115) );
  OAI21_X1 SD1_SB_inst_SD1_SB_bit_inst_40_U29 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_40_n103), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_40_n106), .A(
        SD1_SB_inst_SD1_SB_bit_inst_40_n112), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_40_n113) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_40_U28 ( .A(StateRegOutput[40]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_40_n111), .ZN(OutputRegIn[40]) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_40_U27 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_40_n110), .B2(CipherErrorVec[72]), .A(
        SD1_SB_inst_SD1_SB_bit_inst_40_n109), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_40_n111) );
  AOI221_X1 SD1_SB_inst_SD1_SB_bit_inst_40_U26 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_40_n107), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_40_n112), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_40_n108), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_40_n129), .A(
        SD1_SB_inst_SD1_SB_bit_inst_40_n104), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_40_n109) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_40_U25 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_40_n120), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_40_n112) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_40_U24 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_40_n100), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_40_n102), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_40_n120) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_40_U23 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_40_n130), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_40_n105), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_40_n110) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_40_U22 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_40_n108), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_40_n107) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_40_U21 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_40_n106), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_40_n105) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_40_U20 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_40_n104), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_40_n103) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_40_U19 ( .A(CipherErrorVec[72]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_40_n102) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_40_U18 ( .A(CipherErrorVec[71]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_40_n101) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_40_U17 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_40_n101), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_40_n100) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_40_U16 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_40_n99), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_40_n130) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_40_U15 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_40_n97), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_40_n129) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_40_U14 ( .A(CipherErrorVec[70]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_40_n96) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_40_U13 ( .A(CipherErrorVec[75]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_40_n108) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_40_U12 ( .A(CipherErrorVec[74]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_40_n106) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_40_U11 ( .A(CipherErrorVec[73]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_40_n104) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_40_U10 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_40_n100), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_40_n107), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_40_n98) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_40_U9 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_40_n98), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_40_n104), .A(
        SD1_SB_inst_SD1_SB_bit_inst_40_n96), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_40_n99) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_40_U8 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_40_n105), .A2(CipherErrorVec[72]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_40_n95) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_40_U7 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_40_n95), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_40_n96), .A(
        SD1_SB_inst_SD1_SB_bit_inst_40_n101), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_40_n97) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_40_U6 ( .A(StateRegOutput[41]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_40_n94), .ZN(OutputRegIn[41]) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_40_U5 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_40_n107), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_40_n92), .A(
        SD1_SB_inst_SD1_SB_bit_inst_40_n93), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_40_n94) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_40_U4 ( .A1(CipherErrorVec[72]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_40_n130), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_40_n106), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_40_n93) );
  OAI22_X1 SD1_SB_inst_SD1_SB_bit_inst_40_U3 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_40_n103), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_40_n129), .B1(CipherErrorVec[76]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_40_n128), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_40_n92) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_41_U37 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_41_n110), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_41_n109), .A(
        SD1_SB_inst_SD1_SB_bit_inst_41_n108), .ZN(Feedback[25]) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_41_U36 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_41_n107), .B2(StateRegOutput[40]), .A(
        SD1_SB_inst_SD1_SB_bit_inst_41_n106), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_41_n108) );
  OAI22_X1 SD1_SB_inst_SD1_SB_bit_inst_41_U35 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_41_n109), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_41_n110), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_41_n107), .B2(StateRegOutput[40]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_41_n106) );
  AOI22_X1 SD1_SB_inst_SD1_SB_bit_inst_41_U34 ( .A1(CipherErrorVec[70]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_41_n105), .B1(CipherErrorVec[73]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_41_n104), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_41_n107) );
  OAI21_X1 SD1_SB_inst_SD1_SB_bit_inst_41_U33 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_41_n103), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_41_n102), .A(
        SD1_SB_inst_SD1_SB_bit_inst_41_n101), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_41_n104) );
  NAND3_X1 SD1_SB_inst_SD1_SB_bit_inst_41_U32 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_41_n79), .A2(CipherErrorVec[75]), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_41_n78), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_41_n101) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_41_U31 ( .A1(CipherErrorVec[70]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_41_n79), .A3(CipherErrorVec[74]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_41_n103) );
  AOI211_X1 SD1_SB_inst_SD1_SB_bit_inst_41_U30 ( .C1(
        SD1_SB_inst_SD1_SB_bit_inst_41_n100), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_41_n78), .A(CipherErrorVec[74]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_41_n80), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_41_n105) );
  XOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_41_U29 ( .A(StateRegOutput[42]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_41_n99), .Z(
        SD1_SB_inst_SD1_SB_bit_inst_41_n109) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_41_U28 ( .B1(CipherErrorVec[76]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_41_n98), .A(
        SD1_SB_inst_SD1_SB_bit_inst_41_n97), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_41_n99) );
  AOI221_X1 SD1_SB_inst_SD1_SB_bit_inst_41_U27 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_41_n77), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_41_n96), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_41_n78), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_41_n95), .A(
        SD1_SB_inst_SD1_SB_bit_inst_41_n94), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_41_n97) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_41_U26 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_41_n93), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_41_n94) );
  OAI22_X1 SD1_SB_inst_SD1_SB_bit_inst_41_U25 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_41_n92), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_41_n80), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_41_n91), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_41_n82), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_41_n98) );
  AOI211_X1 SD1_SB_inst_SD1_SB_bit_inst_41_U24 ( .C1(CipherErrorVec[70]), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_41_n100), .A(
        SD1_SB_inst_SD1_SB_bit_inst_41_n79), .B(
        SD1_SB_inst_SD1_SB_bit_inst_41_n90), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_41_n91) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_41_U23 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_41_n102), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_41_n90) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_41_U22 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_41_n77), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_41_n83), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_41_n102) );
  AOI22_X1 SD1_SB_inst_SD1_SB_bit_inst_41_U21 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_41_n77), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_41_n81), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_41_n89), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_41_n83), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_41_n92) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_41_U20 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_41_n77), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_41_n95), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_41_n89) );
  XOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_41_U19 ( .A(StateRegOutput[43]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_41_n88), .Z(
        SD1_SB_inst_SD1_SB_bit_inst_41_n110) );
  OAI21_X1 SD1_SB_inst_SD1_SB_bit_inst_41_U18 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_41_n87), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_41_n96), .A(
        SD1_SB_inst_SD1_SB_bit_inst_41_n86), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_41_n88) );
  OAI221_X1 SD1_SB_inst_SD1_SB_bit_inst_41_U17 ( .B1(CipherErrorVec[74]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_41_n85), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_41_n82), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_41_n84), .A(CipherErrorVec[76]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_41_n86) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_41_U16 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_41_n77), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_41_n79), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_41_n81), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_41_n84) );
  OAI33_X1 SD1_SB_inst_SD1_SB_bit_inst_41_U15 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_41_n79), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_41_n100), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_41_n78), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_41_n80), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_41_n83), .B3(
        SD1_SB_inst_SD1_SB_bit_inst_41_n77), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_41_n85) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_41_U14 ( .A1(CipherErrorVec[73]), .A2(
        CipherErrorVec[75]), .ZN(SD1_SB_inst_SD1_SB_bit_inst_41_n100) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_41_U13 ( .A1(CipherErrorVec[73]), .A2(
        CipherErrorVec[75]), .ZN(SD1_SB_inst_SD1_SB_bit_inst_41_n96) );
  AOI221_X1 SD1_SB_inst_SD1_SB_bit_inst_41_U12 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_41_n93), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_41_n77), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_41_n95), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_41_n77), .A(CipherErrorVec[76]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_41_n87) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_41_U11 ( .A(CipherErrorVec[70]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_41_n95) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_41_U10 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_41_n80), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_41_n82), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_41_n93) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_41_U9 ( .A(CipherErrorVec[73]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_41_n81) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_41_U8 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_41_n80), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_41_n79) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_41_U7 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_41_n78), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_41_n77) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_41_U6 ( .A(CipherErrorVec[74]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_41_n82) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_41_U5 ( .A(CipherErrorVec[75]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_41_n83) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_41_U4 ( .A(CipherErrorVec[72]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_41_n80) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_41_U3 ( .A(CipherErrorVec[71]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_41_n78) );
  OAI22_X1 SD1_SB_inst_SD1_SB_bit_inst_42_U45 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_42_n138), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_42_n137), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_42_n136), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_42_n135), .ZN(Feedback[26]) );
  XOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_42_U44 ( .A(StateRegOutput[41]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_42_n134), .Z(
        SD1_SB_inst_SD1_SB_bit_inst_42_n137) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_42_U43 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_42_n103), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_42_n133), .A(
        SD1_SB_inst_SD1_SB_bit_inst_42_n132), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_42_n134) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_42_U42 ( .A1(CipherErrorVec[73]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_42_n131), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_42_n130), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_42_n132) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_42_U41 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_42_n105), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_42_n99), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_42_n130) );
  OAI22_X1 SD1_SB_inst_SD1_SB_bit_inst_42_U40 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_42_n101), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_42_n129), .B1(CipherErrorVec[76]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_42_n128), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_42_n133) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_42_U39 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_42_n135), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_42_n136), .A(
        SD1_SB_inst_SD1_SB_bit_inst_42_n127), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_42_n138) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_42_U38 ( .A(StateRegOutput[42]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_42_n126), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_42_n127) );
  AOI211_X1 SD1_SB_inst_SD1_SB_bit_inst_42_U37 ( .C1(
        SD1_SB_inst_SD1_SB_bit_inst_42_n101), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_42_n125), .A(
        SD1_SB_inst_SD1_SB_bit_inst_42_n124), .B(
        SD1_SB_inst_SD1_SB_bit_inst_42_n123), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_42_n126) );
  AOI211_X1 SD1_SB_inst_SD1_SB_bit_inst_42_U36 ( .C1(
        SD1_SB_inst_SD1_SB_bit_inst_42_n122), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_42_n102), .A(
        SD1_SB_inst_SD1_SB_bit_inst_42_n121), .B(
        SD1_SB_inst_SD1_SB_bit_inst_42_n104), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_42_n123) );
  AOI22_X1 SD1_SB_inst_SD1_SB_bit_inst_42_U35 ( .A1(CipherErrorVec[70]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_42_n120), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_42_n99), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_42_n106), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_42_n122) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_42_U34 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_42_n102), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_42_n104), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_42_n119), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_42_n124) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_42_U33 ( .A(CipherErrorVec[76]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_42_n121) );
  OAI221_X1 SD1_SB_inst_SD1_SB_bit_inst_42_U32 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_42_n103), .B2(CipherErrorVec[76]), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_42_n103), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_42_n106), .A(CipherErrorVec[70]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_42_n118) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_42_U31 ( .A(StateRegOutput[40]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_42_n117), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_42_n136) );
  AOI22_X1 SD1_SB_inst_SD1_SB_bit_inst_42_U30 ( .A1(CipherErrorVec[73]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_42_n116), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_42_n101), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_42_n115), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_42_n117) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_42_U29 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_42_n103), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_42_n129), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_42_n115) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_42_U28 ( .A1(CipherErrorVec[70]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_42_n114), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_42_n129) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_42_U27 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_42_n120), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_42_n100), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_42_n114) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_42_U26 ( .A1(CipherErrorVec[73]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_42_n105), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_42_n120) );
  OAI21_X1 SD1_SB_inst_SD1_SB_bit_inst_42_U25 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_42_n131), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_42_n113), .A(
        SD1_SB_inst_SD1_SB_bit_inst_42_n128), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_42_n116) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_42_U24 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_42_n99), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_42_n106), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_42_n113) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_42_U23 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_42_n101), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_42_n103), .A3(CipherErrorVec[70]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_42_n131) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_42_U22 ( .A(StateRegOutput[43]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_42_n112), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_42_n135) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_42_U21 ( .B1(CipherErrorVec[76]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_42_n111), .A(
        SD1_SB_inst_SD1_SB_bit_inst_42_n110), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_42_n112) );
  AOI221_X1 SD1_SB_inst_SD1_SB_bit_inst_42_U20 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_42_n104), .B2(CipherErrorVec[70]), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_42_n102), .C2(CipherErrorVec[70]), .A(
        SD1_SB_inst_SD1_SB_bit_inst_42_n119), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_42_n110) );
  NAND3_X1 SD1_SB_inst_SD1_SB_bit_inst_42_U19 ( .A1(CipherErrorVec[73]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_42_n105), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_42_n99), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_42_n119) );
  OAI221_X1 SD1_SB_inst_SD1_SB_bit_inst_42_U18 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_42_n103), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_42_n128), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_42_n103), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_42_n109), .A(
        SD1_SB_inst_SD1_SB_bit_inst_42_n108), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_42_n111) );
  OAI21_X1 SD1_SB_inst_SD1_SB_bit_inst_42_U17 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_42_n105), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_42_n107), .A(CipherErrorVec[73]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_42_n108) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_42_U16 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_42_n101), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_42_n99), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_42_n104), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_42_n107) );
  OAI211_X1 SD1_SB_inst_SD1_SB_bit_inst_42_U15 ( .C1(CipherErrorVec[73]), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_42_n105), .A(
        SD1_SB_inst_SD1_SB_bit_inst_42_n99), .B(
        SD1_SB_inst_SD1_SB_bit_inst_42_n102), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_42_n109) );
  NAND3_X1 SD1_SB_inst_SD1_SB_bit_inst_42_U14 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_42_n101), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_42_n105), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_42_n100), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_42_n128) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_42_U13 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_42_n106), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_42_n105) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_42_U12 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_42_n104), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_42_n103) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_42_U11 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_42_n102), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_42_n101) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_42_U10 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_42_n100), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_42_n99) );
  MUX2_X1 SD1_SB_inst_SD1_SB_bit_inst_42_U9 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_42_n97), .B(
        SD1_SB_inst_SD1_SB_bit_inst_42_n98), .S(
        SD1_SB_inst_SD1_SB_bit_inst_42_n99), .Z(
        SD1_SB_inst_SD1_SB_bit_inst_42_n125) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_42_U8 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_42_n118), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_42_n97) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_42_U7 ( .A(CipherErrorVec[74]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_42_n104) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_42_U6 ( .A(CipherErrorVec[72]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_42_n102) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_42_U5 ( .A(CipherErrorVec[75]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_42_n106) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_42_U4 ( .A(CipherErrorVec[71]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_42_n100) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_42_U3 ( .A1(CipherErrorVec[73]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_42_n121), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_42_n98) );
  AOI222_X1 SD1_SB_inst_SD1_SB_bit_inst_43_U45 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_43_n141), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_43_n140), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_43_n141), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_43_n139), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_43_n140), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_43_n138), .ZN(Feedback[27]) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_43_U44 ( .A(StateRegOutput[40]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_43_n137), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_43_n138) );
  AOI211_X1 SD1_SB_inst_SD1_SB_bit_inst_43_U43 ( .C1(
        SD1_SB_inst_SD1_SB_bit_inst_43_n136), .C2(CipherErrorVec[73]), .A(
        SD1_SB_inst_SD1_SB_bit_inst_43_n135), .B(
        SD1_SB_inst_SD1_SB_bit_inst_43_n134), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_43_n137) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_43_U42 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_43_n105), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_43_n103), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_43_n133), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_43_n134) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_43_U41 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_43_n107), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_43_n132), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_43_n131), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_43_n135) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_43_U40 ( .A1(CipherErrorVec[73]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_43_n100), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_43_n131) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_43_U39 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_43_n130), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_43_n136) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_43_U38 ( .A(StateRegOutput[42]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_43_n129), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_43_n139) );
  AOI22_X1 SD1_SB_inst_SD1_SB_bit_inst_43_U37 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_43_n128), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_43_n127), .B1(CipherErrorVec[76]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_43_n126), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_43_n129) );
  OAI211_X1 SD1_SB_inst_SD1_SB_bit_inst_43_U36 ( .C1(
        SD1_SB_inst_SD1_SB_bit_inst_43_n125), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_43_n101), .A(
        SD1_SB_inst_SD1_SB_bit_inst_43_n124), .B(
        SD1_SB_inst_SD1_SB_bit_inst_43_n123), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_43_n126) );
  NAND3_X1 SD1_SB_inst_SD1_SB_bit_inst_43_U35 ( .A1(CipherErrorVec[70]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_43_n108), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_43_n122), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_43_n123) );
  OAI22_X1 SD1_SB_inst_SD1_SB_bit_inst_43_U34 ( .A1(CipherErrorVec[73]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_43_n106), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_43_n100), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_43_n103), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_43_n122) );
  AOI22_X1 SD1_SB_inst_SD1_SB_bit_inst_43_U33 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_43_n102), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_43_n104), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_43_n105), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_43_n108), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_43_n125) );
  OAI21_X1 SD1_SB_inst_SD1_SB_bit_inst_43_U32 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_43_n100), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_43_n121), .A(
        SD1_SB_inst_SD1_SB_bit_inst_43_n120), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_43_n127) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_43_U31 ( .A(CipherErrorVec[70]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_43_n121) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_43_U30 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_43_n124), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_43_n128) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_43_U29 ( .A(StateRegOutput[41]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_43_n119), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_43_n140) );
  AOI22_X1 SD1_SB_inst_SD1_SB_bit_inst_43_U28 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_43_n105), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_43_n118), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_43_n100), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_43_n117), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_43_n119) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_43_U27 ( .A1(CipherErrorVec[73]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_43_n132), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_43_n108), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_43_n117) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_43_U26 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_43_n102), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_43_n105), .A3(CipherErrorVec[70]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_43_n132) );
  OAI22_X1 SD1_SB_inst_SD1_SB_bit_inst_43_U25 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_43_n102), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_43_n133), .B1(CipherErrorVec[76]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_43_n130), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_43_n118) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_43_U24 ( .A1(CipherErrorVec[70]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_43_n116), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_43_n133) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_43_U23 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_43_n115), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_43_n101), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_43_n116) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_43_U22 ( .A1(CipherErrorVec[73]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_43_n107), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_43_n115) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_43_U21 ( .A(StateRegOutput[43]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_43_n114), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_43_n141) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_43_U20 ( .B1(CipherErrorVec[76]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_43_n113), .A(
        SD1_SB_inst_SD1_SB_bit_inst_43_n112), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_43_n114) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_43_U19 ( .B1(CipherErrorVec[70]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_43_n124), .A(
        SD1_SB_inst_SD1_SB_bit_inst_43_n120), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_43_n112) );
  NAND3_X1 SD1_SB_inst_SD1_SB_bit_inst_43_U18 ( .A1(CipherErrorVec[73]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_43_n100), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_43_n107), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_43_n120) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_43_U17 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_43_n102), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_43_n105), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_43_n124) );
  OAI221_X1 SD1_SB_inst_SD1_SB_bit_inst_43_U16 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_43_n105), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_43_n130), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_43_n105), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_43_n111), .A(
        SD1_SB_inst_SD1_SB_bit_inst_43_n110), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_43_n113) );
  OAI21_X1 SD1_SB_inst_SD1_SB_bit_inst_43_U15 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_43_n107), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_43_n109), .A(CipherErrorVec[73]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_43_n110) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_43_U14 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_43_n102), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_43_n100), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_43_n106), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_43_n109) );
  OAI211_X1 SD1_SB_inst_SD1_SB_bit_inst_43_U13 ( .C1(CipherErrorVec[73]), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_43_n107), .A(
        SD1_SB_inst_SD1_SB_bit_inst_43_n100), .B(
        SD1_SB_inst_SD1_SB_bit_inst_43_n103), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_43_n111) );
  NAND3_X1 SD1_SB_inst_SD1_SB_bit_inst_43_U12 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_43_n102), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_43_n107), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_43_n101), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_43_n130) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_43_U11 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_43_n108), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_43_n107) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_43_U10 ( .A(CipherErrorVec[74]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_43_n106) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_43_U9 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_43_n106), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_43_n105) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_43_U8 ( .A(CipherErrorVec[73]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_43_n104) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_43_U7 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_43_n103), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_43_n102) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_43_U6 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_43_n101), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_43_n100) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_43_U5 ( .A(CipherErrorVec[72]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_43_n103) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_43_U4 ( .A(CipherErrorVec[75]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_43_n108) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_43_U3 ( .A(CipherErrorVec[71]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_43_n101) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_44_U47 ( .B1(OutputRegIn[46]), .B2(
        OutputRegIn[47]), .A(SD1_SB_inst_SD1_SB_bit_inst_44_n131), .ZN(
        Feedback[20]) );
  AOI221_X1 SD1_SB_inst_SD1_SB_bit_inst_44_U46 ( .B1(OutputRegIn[46]), .B2(
        OutputRegIn[44]), .C1(OutputRegIn[47]), .C2(OutputRegIn[44]), .A(
        OutputRegIn[45]), .ZN(SD1_SB_inst_SD1_SB_bit_inst_44_n131) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_44_U45 ( .A(StateRegOutput[47]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_44_n127), .ZN(OutputRegIn[47]) );
  AOI211_X1 SD1_SB_inst_SD1_SB_bit_inst_44_U44 ( .C1(CipherErrorVec[83]), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_44_n126), .A(
        SD1_SB_inst_SD1_SB_bit_inst_44_n125), .B(
        SD1_SB_inst_SD1_SB_bit_inst_44_n124), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_44_n127) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_44_U43 ( .A1(CipherErrorVec[77]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_44_n101), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_44_n123), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_44_n124) );
  AOI222_X1 SD1_SB_inst_SD1_SB_bit_inst_44_U42 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_44_n108), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_44_n104), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_44_n108), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_44_n122), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_44_n104), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_44_n121), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_44_n126) );
  OAI221_X1 SD1_SB_inst_SD1_SB_bit_inst_44_U41 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_44_n120), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_44_n100), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_44_n120), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_44_n102), .A(
        SD1_SB_inst_SD1_SB_bit_inst_44_n106), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_44_n121) );
  OAI211_X1 SD1_SB_inst_SD1_SB_bit_inst_44_U40 ( .C1(
        SD1_SB_inst_SD1_SB_bit_inst_44_n105), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_44_n100), .A(
        SD1_SB_inst_SD1_SB_bit_inst_44_n119), .B(
        SD1_SB_inst_SD1_SB_bit_inst_44_n102), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_44_n122) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_44_U39 ( .A(StateRegOutput[46]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_44_n118), .ZN(OutputRegIn[46]) );
  AOI211_X1 SD1_SB_inst_SD1_SB_bit_inst_44_U38 ( .C1(CipherErrorVec[83]), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_44_n117), .A(
        SD1_SB_inst_SD1_SB_bit_inst_44_n125), .B(
        SD1_SB_inst_SD1_SB_bit_inst_44_n116), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_44_n118) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_44_U37 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_44_n128), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_44_n96), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_44_n116) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_44_U36 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_44_n105), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_44_n120), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_44_n128) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_44_U35 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_44_n102), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_44_n123), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_44_n119), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_44_n125) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_44_U34 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_44_n105), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_44_n100), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_44_n119) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_44_U33 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_44_n107), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_44_n103), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_44_n123) );
  OAI22_X1 SD1_SB_inst_SD1_SB_bit_inst_44_U32 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_44_n107), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_44_n115), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_44_n114), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_44_n102), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_44_n117) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_44_U31 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_44_n100), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_44_n104), .A(
        SD1_SB_inst_SD1_SB_bit_inst_44_n105), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_44_n114) );
  AOI22_X1 SD1_SB_inst_SD1_SB_bit_inst_44_U30 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_44_n105), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_44_n100), .B1(CipherErrorVec[77]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_44_n113), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_44_n115) );
  OAI21_X1 SD1_SB_inst_SD1_SB_bit_inst_44_U29 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_44_n103), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_44_n106), .A(
        SD1_SB_inst_SD1_SB_bit_inst_44_n112), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_44_n113) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_44_U28 ( .A(StateRegOutput[44]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_44_n111), .ZN(OutputRegIn[44]) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_44_U27 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_44_n110), .B2(CipherErrorVec[79]), .A(
        SD1_SB_inst_SD1_SB_bit_inst_44_n109), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_44_n111) );
  AOI221_X1 SD1_SB_inst_SD1_SB_bit_inst_44_U26 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_44_n107), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_44_n112), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_44_n108), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_44_n129), .A(
        SD1_SB_inst_SD1_SB_bit_inst_44_n104), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_44_n109) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_44_U25 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_44_n120), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_44_n112) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_44_U24 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_44_n100), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_44_n102), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_44_n120) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_44_U23 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_44_n130), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_44_n105), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_44_n110) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_44_U22 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_44_n108), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_44_n107) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_44_U21 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_44_n106), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_44_n105) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_44_U20 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_44_n104), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_44_n103) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_44_U19 ( .A(CipherErrorVec[79]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_44_n102) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_44_U18 ( .A(CipherErrorVec[78]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_44_n101) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_44_U17 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_44_n101), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_44_n100) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_44_U16 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_44_n99), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_44_n130) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_44_U15 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_44_n97), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_44_n129) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_44_U14 ( .A(CipherErrorVec[77]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_44_n96) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_44_U13 ( .A(CipherErrorVec[82]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_44_n108) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_44_U12 ( .A(CipherErrorVec[81]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_44_n106) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_44_U11 ( .A(CipherErrorVec[80]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_44_n104) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_44_U10 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_44_n100), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_44_n107), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_44_n98) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_44_U9 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_44_n98), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_44_n104), .A(
        SD1_SB_inst_SD1_SB_bit_inst_44_n96), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_44_n99) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_44_U8 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_44_n105), .A2(CipherErrorVec[79]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_44_n95) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_44_U7 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_44_n95), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_44_n96), .A(
        SD1_SB_inst_SD1_SB_bit_inst_44_n101), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_44_n97) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_44_U6 ( .A(StateRegOutput[45]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_44_n94), .ZN(OutputRegIn[45]) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_44_U5 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_44_n107), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_44_n92), .A(
        SD1_SB_inst_SD1_SB_bit_inst_44_n93), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_44_n94) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_44_U4 ( .A1(CipherErrorVec[79]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_44_n130), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_44_n106), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_44_n93) );
  OAI22_X1 SD1_SB_inst_SD1_SB_bit_inst_44_U3 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_44_n103), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_44_n129), .B1(CipherErrorVec[83]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_44_n128), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_44_n92) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_45_U37 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_45_n110), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_45_n109), .A(
        SD1_SB_inst_SD1_SB_bit_inst_45_n108), .ZN(Feedback[21]) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_45_U36 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_45_n107), .B2(StateRegOutput[44]), .A(
        SD1_SB_inst_SD1_SB_bit_inst_45_n106), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_45_n108) );
  OAI22_X1 SD1_SB_inst_SD1_SB_bit_inst_45_U35 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_45_n109), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_45_n110), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_45_n107), .B2(StateRegOutput[44]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_45_n106) );
  AOI22_X1 SD1_SB_inst_SD1_SB_bit_inst_45_U34 ( .A1(CipherErrorVec[77]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_45_n105), .B1(CipherErrorVec[80]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_45_n104), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_45_n107) );
  OAI21_X1 SD1_SB_inst_SD1_SB_bit_inst_45_U33 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_45_n103), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_45_n102), .A(
        SD1_SB_inst_SD1_SB_bit_inst_45_n101), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_45_n104) );
  NAND3_X1 SD1_SB_inst_SD1_SB_bit_inst_45_U32 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_45_n79), .A2(CipherErrorVec[82]), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_45_n78), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_45_n101) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_45_U31 ( .A1(CipherErrorVec[77]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_45_n79), .A3(CipherErrorVec[81]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_45_n103) );
  AOI211_X1 SD1_SB_inst_SD1_SB_bit_inst_45_U30 ( .C1(
        SD1_SB_inst_SD1_SB_bit_inst_45_n100), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_45_n78), .A(CipherErrorVec[81]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_45_n80), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_45_n105) );
  XOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_45_U29 ( .A(StateRegOutput[46]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_45_n99), .Z(
        SD1_SB_inst_SD1_SB_bit_inst_45_n109) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_45_U28 ( .B1(CipherErrorVec[83]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_45_n98), .A(
        SD1_SB_inst_SD1_SB_bit_inst_45_n97), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_45_n99) );
  AOI221_X1 SD1_SB_inst_SD1_SB_bit_inst_45_U27 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_45_n77), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_45_n96), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_45_n78), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_45_n95), .A(
        SD1_SB_inst_SD1_SB_bit_inst_45_n94), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_45_n97) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_45_U26 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_45_n93), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_45_n94) );
  OAI22_X1 SD1_SB_inst_SD1_SB_bit_inst_45_U25 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_45_n92), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_45_n80), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_45_n91), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_45_n82), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_45_n98) );
  AOI211_X1 SD1_SB_inst_SD1_SB_bit_inst_45_U24 ( .C1(CipherErrorVec[77]), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_45_n100), .A(
        SD1_SB_inst_SD1_SB_bit_inst_45_n79), .B(
        SD1_SB_inst_SD1_SB_bit_inst_45_n90), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_45_n91) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_45_U23 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_45_n102), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_45_n90) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_45_U22 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_45_n77), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_45_n83), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_45_n102) );
  AOI22_X1 SD1_SB_inst_SD1_SB_bit_inst_45_U21 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_45_n77), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_45_n81), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_45_n89), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_45_n83), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_45_n92) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_45_U20 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_45_n77), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_45_n95), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_45_n89) );
  XOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_45_U19 ( .A(StateRegOutput[47]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_45_n88), .Z(
        SD1_SB_inst_SD1_SB_bit_inst_45_n110) );
  OAI21_X1 SD1_SB_inst_SD1_SB_bit_inst_45_U18 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_45_n87), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_45_n96), .A(
        SD1_SB_inst_SD1_SB_bit_inst_45_n86), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_45_n88) );
  OAI221_X1 SD1_SB_inst_SD1_SB_bit_inst_45_U17 ( .B1(CipherErrorVec[81]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_45_n85), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_45_n82), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_45_n84), .A(CipherErrorVec[83]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_45_n86) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_45_U16 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_45_n77), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_45_n79), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_45_n81), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_45_n84) );
  OAI33_X1 SD1_SB_inst_SD1_SB_bit_inst_45_U15 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_45_n79), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_45_n100), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_45_n78), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_45_n80), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_45_n83), .B3(
        SD1_SB_inst_SD1_SB_bit_inst_45_n77), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_45_n85) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_45_U14 ( .A1(CipherErrorVec[80]), .A2(
        CipherErrorVec[82]), .ZN(SD1_SB_inst_SD1_SB_bit_inst_45_n100) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_45_U13 ( .A1(CipherErrorVec[80]), .A2(
        CipherErrorVec[82]), .ZN(SD1_SB_inst_SD1_SB_bit_inst_45_n96) );
  AOI221_X1 SD1_SB_inst_SD1_SB_bit_inst_45_U12 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_45_n93), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_45_n77), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_45_n95), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_45_n77), .A(CipherErrorVec[83]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_45_n87) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_45_U11 ( .A(CipherErrorVec[77]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_45_n95) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_45_U10 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_45_n80), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_45_n82), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_45_n93) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_45_U9 ( .A(CipherErrorVec[80]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_45_n81) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_45_U8 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_45_n80), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_45_n79) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_45_U7 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_45_n78), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_45_n77) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_45_U6 ( .A(CipherErrorVec[81]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_45_n82) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_45_U5 ( .A(CipherErrorVec[82]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_45_n83) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_45_U4 ( .A(CipherErrorVec[79]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_45_n80) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_45_U3 ( .A(CipherErrorVec[78]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_45_n78) );
  OAI22_X1 SD1_SB_inst_SD1_SB_bit_inst_46_U45 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_46_n138), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_46_n137), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_46_n136), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_46_n135), .ZN(Feedback[22]) );
  XOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_46_U44 ( .A(StateRegOutput[45]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_46_n134), .Z(
        SD1_SB_inst_SD1_SB_bit_inst_46_n137) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_46_U43 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_46_n103), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_46_n133), .A(
        SD1_SB_inst_SD1_SB_bit_inst_46_n132), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_46_n134) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_46_U42 ( .A1(CipherErrorVec[80]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_46_n131), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_46_n130), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_46_n132) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_46_U41 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_46_n105), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_46_n99), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_46_n130) );
  OAI22_X1 SD1_SB_inst_SD1_SB_bit_inst_46_U40 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_46_n101), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_46_n129), .B1(CipherErrorVec[83]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_46_n128), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_46_n133) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_46_U39 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_46_n135), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_46_n136), .A(
        SD1_SB_inst_SD1_SB_bit_inst_46_n127), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_46_n138) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_46_U38 ( .A(StateRegOutput[46]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_46_n126), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_46_n127) );
  AOI211_X1 SD1_SB_inst_SD1_SB_bit_inst_46_U37 ( .C1(
        SD1_SB_inst_SD1_SB_bit_inst_46_n101), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_46_n125), .A(
        SD1_SB_inst_SD1_SB_bit_inst_46_n124), .B(
        SD1_SB_inst_SD1_SB_bit_inst_46_n123), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_46_n126) );
  AOI211_X1 SD1_SB_inst_SD1_SB_bit_inst_46_U36 ( .C1(
        SD1_SB_inst_SD1_SB_bit_inst_46_n122), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_46_n102), .A(
        SD1_SB_inst_SD1_SB_bit_inst_46_n121), .B(
        SD1_SB_inst_SD1_SB_bit_inst_46_n104), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_46_n123) );
  AOI22_X1 SD1_SB_inst_SD1_SB_bit_inst_46_U35 ( .A1(CipherErrorVec[77]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_46_n120), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_46_n99), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_46_n106), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_46_n122) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_46_U34 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_46_n102), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_46_n104), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_46_n119), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_46_n124) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_46_U33 ( .A(CipherErrorVec[83]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_46_n121) );
  OAI221_X1 SD1_SB_inst_SD1_SB_bit_inst_46_U32 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_46_n103), .B2(CipherErrorVec[83]), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_46_n103), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_46_n106), .A(CipherErrorVec[77]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_46_n118) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_46_U31 ( .A(StateRegOutput[44]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_46_n117), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_46_n136) );
  AOI22_X1 SD1_SB_inst_SD1_SB_bit_inst_46_U30 ( .A1(CipherErrorVec[80]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_46_n116), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_46_n101), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_46_n115), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_46_n117) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_46_U29 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_46_n103), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_46_n129), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_46_n115) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_46_U28 ( .A1(CipherErrorVec[77]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_46_n114), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_46_n129) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_46_U27 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_46_n120), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_46_n100), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_46_n114) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_46_U26 ( .A1(CipherErrorVec[80]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_46_n105), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_46_n120) );
  OAI21_X1 SD1_SB_inst_SD1_SB_bit_inst_46_U25 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_46_n131), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_46_n113), .A(
        SD1_SB_inst_SD1_SB_bit_inst_46_n128), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_46_n116) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_46_U24 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_46_n99), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_46_n106), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_46_n113) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_46_U23 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_46_n101), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_46_n103), .A3(CipherErrorVec[77]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_46_n131) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_46_U22 ( .A(StateRegOutput[47]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_46_n112), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_46_n135) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_46_U21 ( .B1(CipherErrorVec[83]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_46_n111), .A(
        SD1_SB_inst_SD1_SB_bit_inst_46_n110), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_46_n112) );
  AOI221_X1 SD1_SB_inst_SD1_SB_bit_inst_46_U20 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_46_n104), .B2(CipherErrorVec[77]), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_46_n102), .C2(CipherErrorVec[77]), .A(
        SD1_SB_inst_SD1_SB_bit_inst_46_n119), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_46_n110) );
  NAND3_X1 SD1_SB_inst_SD1_SB_bit_inst_46_U19 ( .A1(CipherErrorVec[80]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_46_n105), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_46_n99), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_46_n119) );
  OAI221_X1 SD1_SB_inst_SD1_SB_bit_inst_46_U18 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_46_n103), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_46_n128), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_46_n103), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_46_n109), .A(
        SD1_SB_inst_SD1_SB_bit_inst_46_n108), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_46_n111) );
  OAI21_X1 SD1_SB_inst_SD1_SB_bit_inst_46_U17 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_46_n105), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_46_n107), .A(CipherErrorVec[80]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_46_n108) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_46_U16 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_46_n101), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_46_n99), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_46_n104), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_46_n107) );
  OAI211_X1 SD1_SB_inst_SD1_SB_bit_inst_46_U15 ( .C1(CipherErrorVec[80]), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_46_n105), .A(
        SD1_SB_inst_SD1_SB_bit_inst_46_n99), .B(
        SD1_SB_inst_SD1_SB_bit_inst_46_n102), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_46_n109) );
  NAND3_X1 SD1_SB_inst_SD1_SB_bit_inst_46_U14 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_46_n101), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_46_n105), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_46_n100), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_46_n128) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_46_U13 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_46_n106), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_46_n105) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_46_U12 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_46_n104), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_46_n103) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_46_U11 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_46_n102), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_46_n101) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_46_U10 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_46_n100), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_46_n99) );
  MUX2_X1 SD1_SB_inst_SD1_SB_bit_inst_46_U9 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_46_n97), .B(
        SD1_SB_inst_SD1_SB_bit_inst_46_n98), .S(
        SD1_SB_inst_SD1_SB_bit_inst_46_n99), .Z(
        SD1_SB_inst_SD1_SB_bit_inst_46_n125) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_46_U8 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_46_n118), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_46_n97) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_46_U7 ( .A(CipherErrorVec[81]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_46_n104) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_46_U6 ( .A(CipherErrorVec[79]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_46_n102) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_46_U5 ( .A(CipherErrorVec[82]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_46_n106) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_46_U4 ( .A(CipherErrorVec[78]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_46_n100) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_46_U3 ( .A1(CipherErrorVec[80]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_46_n121), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_46_n98) );
  AOI222_X1 SD1_SB_inst_SD1_SB_bit_inst_47_U45 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_47_n141), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_47_n140), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_47_n141), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_47_n139), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_47_n140), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_47_n138), .ZN(Feedback[23]) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_47_U44 ( .A(StateRegOutput[44]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_47_n137), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_47_n138) );
  AOI211_X1 SD1_SB_inst_SD1_SB_bit_inst_47_U43 ( .C1(
        SD1_SB_inst_SD1_SB_bit_inst_47_n136), .C2(CipherErrorVec[80]), .A(
        SD1_SB_inst_SD1_SB_bit_inst_47_n135), .B(
        SD1_SB_inst_SD1_SB_bit_inst_47_n134), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_47_n137) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_47_U42 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_47_n105), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_47_n103), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_47_n133), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_47_n134) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_47_U41 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_47_n107), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_47_n132), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_47_n131), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_47_n135) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_47_U40 ( .A1(CipherErrorVec[80]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_47_n100), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_47_n131) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_47_U39 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_47_n130), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_47_n136) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_47_U38 ( .A(StateRegOutput[46]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_47_n129), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_47_n139) );
  AOI22_X1 SD1_SB_inst_SD1_SB_bit_inst_47_U37 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_47_n128), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_47_n127), .B1(CipherErrorVec[83]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_47_n126), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_47_n129) );
  OAI211_X1 SD1_SB_inst_SD1_SB_bit_inst_47_U36 ( .C1(
        SD1_SB_inst_SD1_SB_bit_inst_47_n125), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_47_n101), .A(
        SD1_SB_inst_SD1_SB_bit_inst_47_n124), .B(
        SD1_SB_inst_SD1_SB_bit_inst_47_n123), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_47_n126) );
  NAND3_X1 SD1_SB_inst_SD1_SB_bit_inst_47_U35 ( .A1(CipherErrorVec[77]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_47_n108), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_47_n122), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_47_n123) );
  OAI22_X1 SD1_SB_inst_SD1_SB_bit_inst_47_U34 ( .A1(CipherErrorVec[80]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_47_n106), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_47_n100), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_47_n103), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_47_n122) );
  AOI22_X1 SD1_SB_inst_SD1_SB_bit_inst_47_U33 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_47_n102), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_47_n104), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_47_n105), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_47_n108), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_47_n125) );
  OAI21_X1 SD1_SB_inst_SD1_SB_bit_inst_47_U32 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_47_n100), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_47_n121), .A(
        SD1_SB_inst_SD1_SB_bit_inst_47_n120), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_47_n127) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_47_U31 ( .A(CipherErrorVec[77]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_47_n121) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_47_U30 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_47_n124), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_47_n128) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_47_U29 ( .A(StateRegOutput[45]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_47_n119), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_47_n140) );
  AOI22_X1 SD1_SB_inst_SD1_SB_bit_inst_47_U28 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_47_n105), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_47_n118), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_47_n100), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_47_n117), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_47_n119) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_47_U27 ( .A1(CipherErrorVec[80]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_47_n132), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_47_n108), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_47_n117) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_47_U26 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_47_n102), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_47_n105), .A3(CipherErrorVec[77]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_47_n132) );
  OAI22_X1 SD1_SB_inst_SD1_SB_bit_inst_47_U25 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_47_n102), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_47_n133), .B1(CipherErrorVec[83]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_47_n130), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_47_n118) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_47_U24 ( .A1(CipherErrorVec[77]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_47_n116), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_47_n133) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_47_U23 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_47_n115), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_47_n101), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_47_n116) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_47_U22 ( .A1(CipherErrorVec[80]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_47_n107), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_47_n115) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_47_U21 ( .A(StateRegOutput[47]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_47_n114), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_47_n141) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_47_U20 ( .B1(CipherErrorVec[83]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_47_n113), .A(
        SD1_SB_inst_SD1_SB_bit_inst_47_n112), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_47_n114) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_47_U19 ( .B1(CipherErrorVec[77]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_47_n124), .A(
        SD1_SB_inst_SD1_SB_bit_inst_47_n120), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_47_n112) );
  NAND3_X1 SD1_SB_inst_SD1_SB_bit_inst_47_U18 ( .A1(CipherErrorVec[80]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_47_n100), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_47_n107), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_47_n120) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_47_U17 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_47_n102), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_47_n105), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_47_n124) );
  OAI221_X1 SD1_SB_inst_SD1_SB_bit_inst_47_U16 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_47_n105), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_47_n130), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_47_n105), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_47_n111), .A(
        SD1_SB_inst_SD1_SB_bit_inst_47_n110), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_47_n113) );
  OAI21_X1 SD1_SB_inst_SD1_SB_bit_inst_47_U15 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_47_n107), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_47_n109), .A(CipherErrorVec[80]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_47_n110) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_47_U14 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_47_n102), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_47_n100), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_47_n106), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_47_n109) );
  OAI211_X1 SD1_SB_inst_SD1_SB_bit_inst_47_U13 ( .C1(CipherErrorVec[80]), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_47_n107), .A(
        SD1_SB_inst_SD1_SB_bit_inst_47_n100), .B(
        SD1_SB_inst_SD1_SB_bit_inst_47_n103), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_47_n111) );
  NAND3_X1 SD1_SB_inst_SD1_SB_bit_inst_47_U12 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_47_n102), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_47_n107), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_47_n101), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_47_n130) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_47_U11 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_47_n108), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_47_n107) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_47_U10 ( .A(CipherErrorVec[81]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_47_n106) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_47_U9 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_47_n106), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_47_n105) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_47_U8 ( .A(CipherErrorVec[80]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_47_n104) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_47_U7 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_47_n103), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_47_n102) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_47_U6 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_47_n101), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_47_n100) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_47_U5 ( .A(CipherErrorVec[79]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_47_n103) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_47_U4 ( .A(CipherErrorVec[82]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_47_n108) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_47_U3 ( .A(CipherErrorVec[78]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_47_n101) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_48_U47 ( .B1(OutputRegIn[50]), .B2(
        OutputRegIn[51]), .A(SD1_SB_inst_SD1_SB_bit_inst_48_n131), .ZN(
        Feedback[4]) );
  AOI221_X1 SD1_SB_inst_SD1_SB_bit_inst_48_U46 ( .B1(OutputRegIn[50]), .B2(
        OutputRegIn[48]), .C1(OutputRegIn[51]), .C2(OutputRegIn[48]), .A(
        OutputRegIn[49]), .ZN(SD1_SB_inst_SD1_SB_bit_inst_48_n131) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_48_U45 ( .A(StateRegOutput[51]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_48_n127), .ZN(OutputRegIn[51]) );
  AOI211_X1 SD1_SB_inst_SD1_SB_bit_inst_48_U44 ( .C1(CipherErrorVec[90]), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_48_n126), .A(
        SD1_SB_inst_SD1_SB_bit_inst_48_n125), .B(
        SD1_SB_inst_SD1_SB_bit_inst_48_n124), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_48_n127) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_48_U43 ( .A1(CipherErrorVec[84]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_48_n101), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_48_n123), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_48_n124) );
  AOI222_X1 SD1_SB_inst_SD1_SB_bit_inst_48_U42 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_48_n108), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_48_n104), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_48_n108), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_48_n122), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_48_n104), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_48_n121), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_48_n126) );
  OAI221_X1 SD1_SB_inst_SD1_SB_bit_inst_48_U41 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_48_n120), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_48_n100), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_48_n120), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_48_n102), .A(
        SD1_SB_inst_SD1_SB_bit_inst_48_n106), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_48_n121) );
  OAI211_X1 SD1_SB_inst_SD1_SB_bit_inst_48_U40 ( .C1(
        SD1_SB_inst_SD1_SB_bit_inst_48_n105), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_48_n100), .A(
        SD1_SB_inst_SD1_SB_bit_inst_48_n119), .B(
        SD1_SB_inst_SD1_SB_bit_inst_48_n102), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_48_n122) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_48_U39 ( .A(StateRegOutput[50]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_48_n118), .ZN(OutputRegIn[50]) );
  AOI211_X1 SD1_SB_inst_SD1_SB_bit_inst_48_U38 ( .C1(CipherErrorVec[90]), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_48_n117), .A(
        SD1_SB_inst_SD1_SB_bit_inst_48_n125), .B(
        SD1_SB_inst_SD1_SB_bit_inst_48_n116), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_48_n118) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_48_U37 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_48_n128), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_48_n96), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_48_n116) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_48_U36 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_48_n105), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_48_n120), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_48_n128) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_48_U35 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_48_n102), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_48_n123), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_48_n119), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_48_n125) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_48_U34 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_48_n105), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_48_n100), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_48_n119) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_48_U33 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_48_n107), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_48_n103), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_48_n123) );
  OAI22_X1 SD1_SB_inst_SD1_SB_bit_inst_48_U32 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_48_n107), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_48_n115), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_48_n114), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_48_n102), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_48_n117) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_48_U31 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_48_n100), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_48_n104), .A(
        SD1_SB_inst_SD1_SB_bit_inst_48_n105), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_48_n114) );
  AOI22_X1 SD1_SB_inst_SD1_SB_bit_inst_48_U30 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_48_n105), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_48_n100), .B1(CipherErrorVec[84]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_48_n113), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_48_n115) );
  OAI21_X1 SD1_SB_inst_SD1_SB_bit_inst_48_U29 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_48_n103), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_48_n106), .A(
        SD1_SB_inst_SD1_SB_bit_inst_48_n112), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_48_n113) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_48_U28 ( .A(StateRegOutput[48]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_48_n111), .ZN(OutputRegIn[48]) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_48_U27 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_48_n110), .B2(CipherErrorVec[86]), .A(
        SD1_SB_inst_SD1_SB_bit_inst_48_n109), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_48_n111) );
  AOI221_X1 SD1_SB_inst_SD1_SB_bit_inst_48_U26 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_48_n107), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_48_n112), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_48_n108), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_48_n129), .A(
        SD1_SB_inst_SD1_SB_bit_inst_48_n104), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_48_n109) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_48_U25 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_48_n120), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_48_n112) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_48_U24 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_48_n100), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_48_n102), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_48_n120) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_48_U23 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_48_n130), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_48_n105), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_48_n110) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_48_U22 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_48_n108), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_48_n107) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_48_U21 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_48_n106), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_48_n105) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_48_U20 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_48_n104), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_48_n103) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_48_U19 ( .A(CipherErrorVec[86]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_48_n102) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_48_U18 ( .A(CipherErrorVec[85]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_48_n101) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_48_U17 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_48_n101), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_48_n100) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_48_U16 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_48_n99), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_48_n130) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_48_U15 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_48_n97), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_48_n129) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_48_U14 ( .A(CipherErrorVec[84]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_48_n96) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_48_U13 ( .A(CipherErrorVec[89]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_48_n108) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_48_U12 ( .A(CipherErrorVec[88]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_48_n106) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_48_U11 ( .A(CipherErrorVec[87]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_48_n104) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_48_U10 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_48_n100), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_48_n107), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_48_n98) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_48_U9 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_48_n98), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_48_n104), .A(
        SD1_SB_inst_SD1_SB_bit_inst_48_n96), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_48_n99) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_48_U8 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_48_n105), .A2(CipherErrorVec[86]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_48_n95) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_48_U7 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_48_n95), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_48_n96), .A(
        SD1_SB_inst_SD1_SB_bit_inst_48_n101), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_48_n97) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_48_U6 ( .A(StateRegOutput[49]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_48_n94), .ZN(OutputRegIn[49]) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_48_U5 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_48_n107), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_48_n92), .A(
        SD1_SB_inst_SD1_SB_bit_inst_48_n93), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_48_n94) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_48_U4 ( .A1(CipherErrorVec[86]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_48_n130), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_48_n106), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_48_n93) );
  OAI22_X1 SD1_SB_inst_SD1_SB_bit_inst_48_U3 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_48_n103), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_48_n129), .B1(CipherErrorVec[90]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_48_n128), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_48_n92) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_49_U37 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_49_n110), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_49_n109), .A(
        SD1_SB_inst_SD1_SB_bit_inst_49_n108), .ZN(Feedback[5]) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_49_U36 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_49_n107), .B2(StateRegOutput[48]), .A(
        SD1_SB_inst_SD1_SB_bit_inst_49_n106), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_49_n108) );
  OAI22_X1 SD1_SB_inst_SD1_SB_bit_inst_49_U35 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_49_n109), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_49_n110), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_49_n107), .B2(StateRegOutput[48]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_49_n106) );
  AOI22_X1 SD1_SB_inst_SD1_SB_bit_inst_49_U34 ( .A1(CipherErrorVec[84]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_49_n105), .B1(CipherErrorVec[87]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_49_n104), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_49_n107) );
  OAI21_X1 SD1_SB_inst_SD1_SB_bit_inst_49_U33 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_49_n103), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_49_n102), .A(
        SD1_SB_inst_SD1_SB_bit_inst_49_n101), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_49_n104) );
  NAND3_X1 SD1_SB_inst_SD1_SB_bit_inst_49_U32 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_49_n79), .A2(CipherErrorVec[89]), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_49_n78), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_49_n101) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_49_U31 ( .A1(CipherErrorVec[84]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_49_n79), .A3(CipherErrorVec[88]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_49_n103) );
  AOI211_X1 SD1_SB_inst_SD1_SB_bit_inst_49_U30 ( .C1(
        SD1_SB_inst_SD1_SB_bit_inst_49_n100), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_49_n78), .A(CipherErrorVec[88]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_49_n80), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_49_n105) );
  XOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_49_U29 ( .A(StateRegOutput[50]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_49_n99), .Z(
        SD1_SB_inst_SD1_SB_bit_inst_49_n109) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_49_U28 ( .B1(CipherErrorVec[90]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_49_n98), .A(
        SD1_SB_inst_SD1_SB_bit_inst_49_n97), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_49_n99) );
  AOI221_X1 SD1_SB_inst_SD1_SB_bit_inst_49_U27 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_49_n77), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_49_n96), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_49_n78), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_49_n95), .A(
        SD1_SB_inst_SD1_SB_bit_inst_49_n94), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_49_n97) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_49_U26 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_49_n93), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_49_n94) );
  OAI22_X1 SD1_SB_inst_SD1_SB_bit_inst_49_U25 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_49_n92), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_49_n80), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_49_n91), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_49_n82), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_49_n98) );
  AOI211_X1 SD1_SB_inst_SD1_SB_bit_inst_49_U24 ( .C1(CipherErrorVec[84]), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_49_n100), .A(
        SD1_SB_inst_SD1_SB_bit_inst_49_n79), .B(
        SD1_SB_inst_SD1_SB_bit_inst_49_n90), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_49_n91) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_49_U23 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_49_n102), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_49_n90) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_49_U22 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_49_n77), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_49_n83), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_49_n102) );
  AOI22_X1 SD1_SB_inst_SD1_SB_bit_inst_49_U21 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_49_n77), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_49_n81), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_49_n89), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_49_n83), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_49_n92) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_49_U20 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_49_n77), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_49_n95), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_49_n89) );
  XOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_49_U19 ( .A(StateRegOutput[51]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_49_n88), .Z(
        SD1_SB_inst_SD1_SB_bit_inst_49_n110) );
  OAI21_X1 SD1_SB_inst_SD1_SB_bit_inst_49_U18 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_49_n87), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_49_n96), .A(
        SD1_SB_inst_SD1_SB_bit_inst_49_n86), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_49_n88) );
  OAI221_X1 SD1_SB_inst_SD1_SB_bit_inst_49_U17 ( .B1(CipherErrorVec[88]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_49_n85), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_49_n82), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_49_n84), .A(CipherErrorVec[90]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_49_n86) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_49_U16 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_49_n77), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_49_n79), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_49_n81), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_49_n84) );
  OAI33_X1 SD1_SB_inst_SD1_SB_bit_inst_49_U15 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_49_n79), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_49_n100), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_49_n78), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_49_n80), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_49_n83), .B3(
        SD1_SB_inst_SD1_SB_bit_inst_49_n77), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_49_n85) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_49_U14 ( .A1(CipherErrorVec[87]), .A2(
        CipherErrorVec[89]), .ZN(SD1_SB_inst_SD1_SB_bit_inst_49_n100) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_49_U13 ( .A1(CipherErrorVec[87]), .A2(
        CipherErrorVec[89]), .ZN(SD1_SB_inst_SD1_SB_bit_inst_49_n96) );
  AOI221_X1 SD1_SB_inst_SD1_SB_bit_inst_49_U12 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_49_n93), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_49_n77), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_49_n95), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_49_n77), .A(CipherErrorVec[90]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_49_n87) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_49_U11 ( .A(CipherErrorVec[84]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_49_n95) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_49_U10 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_49_n80), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_49_n82), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_49_n93) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_49_U9 ( .A(CipherErrorVec[87]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_49_n81) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_49_U8 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_49_n80), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_49_n79) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_49_U7 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_49_n78), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_49_n77) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_49_U6 ( .A(CipherErrorVec[88]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_49_n82) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_49_U5 ( .A(CipherErrorVec[89]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_49_n83) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_49_U4 ( .A(CipherErrorVec[86]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_49_n80) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_49_U3 ( .A(CipherErrorVec[85]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_49_n78) );
  OAI22_X1 SD1_SB_inst_SD1_SB_bit_inst_50_U45 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_50_n138), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_50_n137), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_50_n136), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_50_n135), .ZN(Feedback[6]) );
  XOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_50_U44 ( .A(StateRegOutput[49]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_50_n134), .Z(
        SD1_SB_inst_SD1_SB_bit_inst_50_n137) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_50_U43 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_50_n103), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_50_n133), .A(
        SD1_SB_inst_SD1_SB_bit_inst_50_n132), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_50_n134) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_50_U42 ( .A1(CipherErrorVec[87]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_50_n131), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_50_n130), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_50_n132) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_50_U41 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_50_n105), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_50_n99), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_50_n130) );
  OAI22_X1 SD1_SB_inst_SD1_SB_bit_inst_50_U40 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_50_n101), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_50_n129), .B1(CipherErrorVec[90]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_50_n128), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_50_n133) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_50_U39 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_50_n135), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_50_n136), .A(
        SD1_SB_inst_SD1_SB_bit_inst_50_n127), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_50_n138) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_50_U38 ( .A(StateRegOutput[50]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_50_n126), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_50_n127) );
  AOI211_X1 SD1_SB_inst_SD1_SB_bit_inst_50_U37 ( .C1(
        SD1_SB_inst_SD1_SB_bit_inst_50_n101), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_50_n125), .A(
        SD1_SB_inst_SD1_SB_bit_inst_50_n124), .B(
        SD1_SB_inst_SD1_SB_bit_inst_50_n123), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_50_n126) );
  AOI211_X1 SD1_SB_inst_SD1_SB_bit_inst_50_U36 ( .C1(
        SD1_SB_inst_SD1_SB_bit_inst_50_n122), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_50_n102), .A(
        SD1_SB_inst_SD1_SB_bit_inst_50_n121), .B(
        SD1_SB_inst_SD1_SB_bit_inst_50_n104), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_50_n123) );
  AOI22_X1 SD1_SB_inst_SD1_SB_bit_inst_50_U35 ( .A1(CipherErrorVec[84]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_50_n120), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_50_n99), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_50_n106), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_50_n122) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_50_U34 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_50_n102), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_50_n104), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_50_n119), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_50_n124) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_50_U33 ( .A(CipherErrorVec[90]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_50_n121) );
  OAI221_X1 SD1_SB_inst_SD1_SB_bit_inst_50_U32 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_50_n103), .B2(CipherErrorVec[90]), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_50_n103), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_50_n106), .A(CipherErrorVec[84]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_50_n118) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_50_U31 ( .A(StateRegOutput[48]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_50_n117), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_50_n136) );
  AOI22_X1 SD1_SB_inst_SD1_SB_bit_inst_50_U30 ( .A1(CipherErrorVec[87]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_50_n116), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_50_n101), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_50_n115), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_50_n117) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_50_U29 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_50_n103), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_50_n129), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_50_n115) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_50_U28 ( .A1(CipherErrorVec[84]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_50_n114), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_50_n129) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_50_U27 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_50_n120), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_50_n100), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_50_n114) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_50_U26 ( .A1(CipherErrorVec[87]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_50_n105), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_50_n120) );
  OAI21_X1 SD1_SB_inst_SD1_SB_bit_inst_50_U25 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_50_n131), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_50_n113), .A(
        SD1_SB_inst_SD1_SB_bit_inst_50_n128), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_50_n116) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_50_U24 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_50_n99), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_50_n106), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_50_n113) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_50_U23 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_50_n101), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_50_n103), .A3(CipherErrorVec[84]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_50_n131) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_50_U22 ( .A(StateRegOutput[51]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_50_n112), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_50_n135) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_50_U21 ( .B1(CipherErrorVec[90]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_50_n111), .A(
        SD1_SB_inst_SD1_SB_bit_inst_50_n110), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_50_n112) );
  AOI221_X1 SD1_SB_inst_SD1_SB_bit_inst_50_U20 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_50_n104), .B2(CipherErrorVec[84]), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_50_n102), .C2(CipherErrorVec[84]), .A(
        SD1_SB_inst_SD1_SB_bit_inst_50_n119), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_50_n110) );
  NAND3_X1 SD1_SB_inst_SD1_SB_bit_inst_50_U19 ( .A1(CipherErrorVec[87]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_50_n105), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_50_n99), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_50_n119) );
  OAI221_X1 SD1_SB_inst_SD1_SB_bit_inst_50_U18 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_50_n103), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_50_n128), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_50_n103), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_50_n109), .A(
        SD1_SB_inst_SD1_SB_bit_inst_50_n108), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_50_n111) );
  OAI21_X1 SD1_SB_inst_SD1_SB_bit_inst_50_U17 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_50_n105), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_50_n107), .A(CipherErrorVec[87]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_50_n108) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_50_U16 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_50_n101), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_50_n99), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_50_n104), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_50_n107) );
  OAI211_X1 SD1_SB_inst_SD1_SB_bit_inst_50_U15 ( .C1(CipherErrorVec[87]), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_50_n105), .A(
        SD1_SB_inst_SD1_SB_bit_inst_50_n99), .B(
        SD1_SB_inst_SD1_SB_bit_inst_50_n102), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_50_n109) );
  NAND3_X1 SD1_SB_inst_SD1_SB_bit_inst_50_U14 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_50_n101), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_50_n105), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_50_n100), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_50_n128) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_50_U13 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_50_n106), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_50_n105) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_50_U12 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_50_n104), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_50_n103) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_50_U11 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_50_n102), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_50_n101) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_50_U10 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_50_n100), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_50_n99) );
  MUX2_X1 SD1_SB_inst_SD1_SB_bit_inst_50_U9 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_50_n97), .B(
        SD1_SB_inst_SD1_SB_bit_inst_50_n98), .S(
        SD1_SB_inst_SD1_SB_bit_inst_50_n99), .Z(
        SD1_SB_inst_SD1_SB_bit_inst_50_n125) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_50_U8 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_50_n118), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_50_n97) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_50_U7 ( .A(CipherErrorVec[88]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_50_n104) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_50_U6 ( .A(CipherErrorVec[86]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_50_n102) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_50_U5 ( .A(CipherErrorVec[89]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_50_n106) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_50_U4 ( .A(CipherErrorVec[85]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_50_n100) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_50_U3 ( .A1(CipherErrorVec[87]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_50_n121), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_50_n98) );
  AOI222_X1 SD1_SB_inst_SD1_SB_bit_inst_51_U45 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_51_n141), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_51_n140), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_51_n141), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_51_n139), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_51_n140), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_51_n138), .ZN(Feedback[7]) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_51_U44 ( .A(StateRegOutput[48]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_51_n137), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_51_n138) );
  AOI211_X1 SD1_SB_inst_SD1_SB_bit_inst_51_U43 ( .C1(
        SD1_SB_inst_SD1_SB_bit_inst_51_n136), .C2(CipherErrorVec[87]), .A(
        SD1_SB_inst_SD1_SB_bit_inst_51_n135), .B(
        SD1_SB_inst_SD1_SB_bit_inst_51_n134), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_51_n137) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_51_U42 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_51_n105), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_51_n103), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_51_n133), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_51_n134) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_51_U41 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_51_n107), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_51_n132), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_51_n131), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_51_n135) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_51_U40 ( .A1(CipherErrorVec[87]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_51_n100), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_51_n131) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_51_U39 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_51_n130), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_51_n136) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_51_U38 ( .A(StateRegOutput[50]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_51_n129), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_51_n139) );
  AOI22_X1 SD1_SB_inst_SD1_SB_bit_inst_51_U37 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_51_n128), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_51_n127), .B1(CipherErrorVec[90]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_51_n126), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_51_n129) );
  OAI211_X1 SD1_SB_inst_SD1_SB_bit_inst_51_U36 ( .C1(
        SD1_SB_inst_SD1_SB_bit_inst_51_n125), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_51_n101), .A(
        SD1_SB_inst_SD1_SB_bit_inst_51_n124), .B(
        SD1_SB_inst_SD1_SB_bit_inst_51_n123), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_51_n126) );
  NAND3_X1 SD1_SB_inst_SD1_SB_bit_inst_51_U35 ( .A1(CipherErrorVec[84]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_51_n108), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_51_n122), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_51_n123) );
  OAI22_X1 SD1_SB_inst_SD1_SB_bit_inst_51_U34 ( .A1(CipherErrorVec[87]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_51_n106), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_51_n100), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_51_n103), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_51_n122) );
  AOI22_X1 SD1_SB_inst_SD1_SB_bit_inst_51_U33 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_51_n102), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_51_n104), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_51_n105), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_51_n108), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_51_n125) );
  OAI21_X1 SD1_SB_inst_SD1_SB_bit_inst_51_U32 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_51_n100), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_51_n121), .A(
        SD1_SB_inst_SD1_SB_bit_inst_51_n120), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_51_n127) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_51_U31 ( .A(CipherErrorVec[84]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_51_n121) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_51_U30 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_51_n124), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_51_n128) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_51_U29 ( .A(StateRegOutput[49]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_51_n119), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_51_n140) );
  AOI22_X1 SD1_SB_inst_SD1_SB_bit_inst_51_U28 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_51_n105), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_51_n118), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_51_n100), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_51_n117), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_51_n119) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_51_U27 ( .A1(CipherErrorVec[87]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_51_n132), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_51_n108), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_51_n117) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_51_U26 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_51_n102), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_51_n105), .A3(CipherErrorVec[84]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_51_n132) );
  OAI22_X1 SD1_SB_inst_SD1_SB_bit_inst_51_U25 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_51_n102), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_51_n133), .B1(CipherErrorVec[90]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_51_n130), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_51_n118) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_51_U24 ( .A1(CipherErrorVec[84]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_51_n116), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_51_n133) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_51_U23 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_51_n115), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_51_n101), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_51_n116) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_51_U22 ( .A1(CipherErrorVec[87]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_51_n107), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_51_n115) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_51_U21 ( .A(StateRegOutput[51]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_51_n114), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_51_n141) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_51_U20 ( .B1(CipherErrorVec[90]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_51_n113), .A(
        SD1_SB_inst_SD1_SB_bit_inst_51_n112), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_51_n114) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_51_U19 ( .B1(CipherErrorVec[84]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_51_n124), .A(
        SD1_SB_inst_SD1_SB_bit_inst_51_n120), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_51_n112) );
  NAND3_X1 SD1_SB_inst_SD1_SB_bit_inst_51_U18 ( .A1(CipherErrorVec[87]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_51_n100), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_51_n107), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_51_n120) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_51_U17 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_51_n102), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_51_n105), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_51_n124) );
  OAI221_X1 SD1_SB_inst_SD1_SB_bit_inst_51_U16 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_51_n105), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_51_n130), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_51_n105), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_51_n111), .A(
        SD1_SB_inst_SD1_SB_bit_inst_51_n110), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_51_n113) );
  OAI21_X1 SD1_SB_inst_SD1_SB_bit_inst_51_U15 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_51_n107), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_51_n109), .A(CipherErrorVec[87]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_51_n110) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_51_U14 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_51_n102), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_51_n100), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_51_n106), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_51_n109) );
  OAI211_X1 SD1_SB_inst_SD1_SB_bit_inst_51_U13 ( .C1(CipherErrorVec[87]), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_51_n107), .A(
        SD1_SB_inst_SD1_SB_bit_inst_51_n100), .B(
        SD1_SB_inst_SD1_SB_bit_inst_51_n103), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_51_n111) );
  NAND3_X1 SD1_SB_inst_SD1_SB_bit_inst_51_U12 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_51_n102), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_51_n107), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_51_n101), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_51_n130) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_51_U11 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_51_n108), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_51_n107) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_51_U10 ( .A(CipherErrorVec[88]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_51_n106) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_51_U9 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_51_n106), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_51_n105) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_51_U8 ( .A(CipherErrorVec[87]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_51_n104) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_51_U7 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_51_n103), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_51_n102) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_51_U6 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_51_n101), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_51_n100) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_51_U5 ( .A(CipherErrorVec[86]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_51_n103) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_51_U4 ( .A(CipherErrorVec[89]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_51_n108) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_51_U3 ( .A(CipherErrorVec[85]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_51_n101) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_52_U47 ( .B1(OutputRegIn[54]), .B2(
        OutputRegIn[55]), .A(SD1_SB_inst_SD1_SB_bit_inst_52_n131), .ZN(
        Feedback[8]) );
  AOI221_X1 SD1_SB_inst_SD1_SB_bit_inst_52_U46 ( .B1(OutputRegIn[54]), .B2(
        OutputRegIn[52]), .C1(OutputRegIn[55]), .C2(OutputRegIn[52]), .A(
        OutputRegIn[53]), .ZN(SD1_SB_inst_SD1_SB_bit_inst_52_n131) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_52_U45 ( .A(StateRegOutput[55]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_52_n127), .ZN(OutputRegIn[55]) );
  AOI211_X1 SD1_SB_inst_SD1_SB_bit_inst_52_U44 ( .C1(CipherErrorVec[97]), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_52_n126), .A(
        SD1_SB_inst_SD1_SB_bit_inst_52_n125), .B(
        SD1_SB_inst_SD1_SB_bit_inst_52_n124), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_52_n127) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_52_U43 ( .A1(CipherErrorVec[91]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_52_n101), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_52_n123), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_52_n124) );
  AOI222_X1 SD1_SB_inst_SD1_SB_bit_inst_52_U42 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_52_n108), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_52_n104), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_52_n108), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_52_n122), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_52_n104), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_52_n121), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_52_n126) );
  OAI221_X1 SD1_SB_inst_SD1_SB_bit_inst_52_U41 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_52_n120), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_52_n100), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_52_n120), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_52_n102), .A(
        SD1_SB_inst_SD1_SB_bit_inst_52_n106), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_52_n121) );
  OAI211_X1 SD1_SB_inst_SD1_SB_bit_inst_52_U40 ( .C1(
        SD1_SB_inst_SD1_SB_bit_inst_52_n105), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_52_n100), .A(
        SD1_SB_inst_SD1_SB_bit_inst_52_n119), .B(
        SD1_SB_inst_SD1_SB_bit_inst_52_n102), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_52_n122) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_52_U39 ( .A(StateRegOutput[54]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_52_n118), .ZN(OutputRegIn[54]) );
  AOI211_X1 SD1_SB_inst_SD1_SB_bit_inst_52_U38 ( .C1(CipherErrorVec[97]), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_52_n117), .A(
        SD1_SB_inst_SD1_SB_bit_inst_52_n125), .B(
        SD1_SB_inst_SD1_SB_bit_inst_52_n116), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_52_n118) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_52_U37 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_52_n128), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_52_n96), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_52_n116) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_52_U36 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_52_n105), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_52_n120), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_52_n128) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_52_U35 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_52_n102), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_52_n123), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_52_n119), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_52_n125) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_52_U34 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_52_n105), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_52_n100), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_52_n119) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_52_U33 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_52_n107), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_52_n103), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_52_n123) );
  OAI22_X1 SD1_SB_inst_SD1_SB_bit_inst_52_U32 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_52_n107), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_52_n115), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_52_n114), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_52_n102), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_52_n117) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_52_U31 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_52_n100), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_52_n104), .A(
        SD1_SB_inst_SD1_SB_bit_inst_52_n105), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_52_n114) );
  AOI22_X1 SD1_SB_inst_SD1_SB_bit_inst_52_U30 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_52_n105), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_52_n100), .B1(CipherErrorVec[91]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_52_n113), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_52_n115) );
  OAI21_X1 SD1_SB_inst_SD1_SB_bit_inst_52_U29 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_52_n103), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_52_n106), .A(
        SD1_SB_inst_SD1_SB_bit_inst_52_n112), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_52_n113) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_52_U28 ( .A(StateRegOutput[52]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_52_n111), .ZN(OutputRegIn[52]) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_52_U27 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_52_n110), .B2(CipherErrorVec[93]), .A(
        SD1_SB_inst_SD1_SB_bit_inst_52_n109), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_52_n111) );
  AOI221_X1 SD1_SB_inst_SD1_SB_bit_inst_52_U26 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_52_n107), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_52_n112), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_52_n108), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_52_n129), .A(
        SD1_SB_inst_SD1_SB_bit_inst_52_n104), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_52_n109) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_52_U25 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_52_n120), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_52_n112) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_52_U24 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_52_n100), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_52_n102), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_52_n120) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_52_U23 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_52_n130), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_52_n105), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_52_n110) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_52_U22 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_52_n108), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_52_n107) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_52_U21 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_52_n106), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_52_n105) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_52_U20 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_52_n104), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_52_n103) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_52_U19 ( .A(CipherErrorVec[93]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_52_n102) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_52_U18 ( .A(CipherErrorVec[92]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_52_n101) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_52_U17 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_52_n101), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_52_n100) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_52_U16 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_52_n99), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_52_n130) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_52_U15 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_52_n97), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_52_n129) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_52_U14 ( .A(CipherErrorVec[91]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_52_n96) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_52_U13 ( .A(CipherErrorVec[96]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_52_n108) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_52_U12 ( .A(CipherErrorVec[95]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_52_n106) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_52_U11 ( .A(CipherErrorVec[94]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_52_n104) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_52_U10 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_52_n100), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_52_n107), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_52_n98) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_52_U9 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_52_n98), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_52_n104), .A(
        SD1_SB_inst_SD1_SB_bit_inst_52_n96), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_52_n99) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_52_U8 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_52_n105), .A2(CipherErrorVec[93]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_52_n95) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_52_U7 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_52_n95), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_52_n96), .A(
        SD1_SB_inst_SD1_SB_bit_inst_52_n101), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_52_n97) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_52_U6 ( .A(StateRegOutput[53]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_52_n94), .ZN(OutputRegIn[53]) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_52_U5 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_52_n107), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_52_n92), .A(
        SD1_SB_inst_SD1_SB_bit_inst_52_n93), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_52_n94) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_52_U4 ( .A1(CipherErrorVec[93]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_52_n130), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_52_n106), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_52_n93) );
  OAI22_X1 SD1_SB_inst_SD1_SB_bit_inst_52_U3 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_52_n103), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_52_n129), .B1(CipherErrorVec[97]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_52_n128), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_52_n92) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_53_U37 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_53_n110), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_53_n109), .A(
        SD1_SB_inst_SD1_SB_bit_inst_53_n108), .ZN(Feedback[9]) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_53_U36 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_53_n107), .B2(StateRegOutput[52]), .A(
        SD1_SB_inst_SD1_SB_bit_inst_53_n106), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_53_n108) );
  OAI22_X1 SD1_SB_inst_SD1_SB_bit_inst_53_U35 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_53_n109), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_53_n110), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_53_n107), .B2(StateRegOutput[52]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_53_n106) );
  AOI22_X1 SD1_SB_inst_SD1_SB_bit_inst_53_U34 ( .A1(CipherErrorVec[91]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_53_n105), .B1(CipherErrorVec[94]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_53_n104), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_53_n107) );
  OAI21_X1 SD1_SB_inst_SD1_SB_bit_inst_53_U33 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_53_n103), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_53_n102), .A(
        SD1_SB_inst_SD1_SB_bit_inst_53_n101), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_53_n104) );
  NAND3_X1 SD1_SB_inst_SD1_SB_bit_inst_53_U32 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_53_n79), .A2(CipherErrorVec[96]), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_53_n78), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_53_n101) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_53_U31 ( .A1(CipherErrorVec[91]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_53_n79), .A3(CipherErrorVec[95]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_53_n103) );
  AOI211_X1 SD1_SB_inst_SD1_SB_bit_inst_53_U30 ( .C1(
        SD1_SB_inst_SD1_SB_bit_inst_53_n100), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_53_n78), .A(CipherErrorVec[95]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_53_n80), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_53_n105) );
  XOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_53_U29 ( .A(StateRegOutput[54]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_53_n99), .Z(
        SD1_SB_inst_SD1_SB_bit_inst_53_n109) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_53_U28 ( .B1(CipherErrorVec[97]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_53_n98), .A(
        SD1_SB_inst_SD1_SB_bit_inst_53_n97), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_53_n99) );
  AOI221_X1 SD1_SB_inst_SD1_SB_bit_inst_53_U27 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_53_n77), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_53_n96), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_53_n78), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_53_n95), .A(
        SD1_SB_inst_SD1_SB_bit_inst_53_n94), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_53_n97) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_53_U26 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_53_n93), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_53_n94) );
  OAI22_X1 SD1_SB_inst_SD1_SB_bit_inst_53_U25 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_53_n92), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_53_n80), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_53_n91), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_53_n82), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_53_n98) );
  AOI211_X1 SD1_SB_inst_SD1_SB_bit_inst_53_U24 ( .C1(CipherErrorVec[91]), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_53_n100), .A(
        SD1_SB_inst_SD1_SB_bit_inst_53_n79), .B(
        SD1_SB_inst_SD1_SB_bit_inst_53_n90), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_53_n91) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_53_U23 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_53_n102), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_53_n90) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_53_U22 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_53_n77), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_53_n83), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_53_n102) );
  AOI22_X1 SD1_SB_inst_SD1_SB_bit_inst_53_U21 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_53_n77), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_53_n81), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_53_n89), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_53_n83), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_53_n92) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_53_U20 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_53_n77), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_53_n95), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_53_n89) );
  XOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_53_U19 ( .A(StateRegOutput[55]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_53_n88), .Z(
        SD1_SB_inst_SD1_SB_bit_inst_53_n110) );
  OAI21_X1 SD1_SB_inst_SD1_SB_bit_inst_53_U18 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_53_n87), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_53_n96), .A(
        SD1_SB_inst_SD1_SB_bit_inst_53_n86), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_53_n88) );
  OAI221_X1 SD1_SB_inst_SD1_SB_bit_inst_53_U17 ( .B1(CipherErrorVec[95]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_53_n85), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_53_n82), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_53_n84), .A(CipherErrorVec[97]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_53_n86) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_53_U16 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_53_n77), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_53_n79), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_53_n81), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_53_n84) );
  OAI33_X1 SD1_SB_inst_SD1_SB_bit_inst_53_U15 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_53_n79), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_53_n100), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_53_n78), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_53_n80), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_53_n83), .B3(
        SD1_SB_inst_SD1_SB_bit_inst_53_n77), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_53_n85) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_53_U14 ( .A1(CipherErrorVec[94]), .A2(
        CipherErrorVec[96]), .ZN(SD1_SB_inst_SD1_SB_bit_inst_53_n100) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_53_U13 ( .A1(CipherErrorVec[94]), .A2(
        CipherErrorVec[96]), .ZN(SD1_SB_inst_SD1_SB_bit_inst_53_n96) );
  AOI221_X1 SD1_SB_inst_SD1_SB_bit_inst_53_U12 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_53_n93), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_53_n77), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_53_n95), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_53_n77), .A(CipherErrorVec[97]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_53_n87) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_53_U11 ( .A(CipherErrorVec[91]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_53_n95) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_53_U10 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_53_n80), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_53_n82), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_53_n93) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_53_U9 ( .A(CipherErrorVec[94]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_53_n81) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_53_U8 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_53_n80), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_53_n79) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_53_U7 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_53_n78), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_53_n77) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_53_U6 ( .A(CipherErrorVec[95]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_53_n82) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_53_U5 ( .A(CipherErrorVec[96]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_53_n83) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_53_U4 ( .A(CipherErrorVec[93]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_53_n80) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_53_U3 ( .A(CipherErrorVec[92]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_53_n78) );
  OAI22_X1 SD1_SB_inst_SD1_SB_bit_inst_54_U45 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_54_n138), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_54_n137), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_54_n136), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_54_n135), .ZN(Feedback[10]) );
  XOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_54_U44 ( .A(StateRegOutput[53]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_54_n134), .Z(
        SD1_SB_inst_SD1_SB_bit_inst_54_n137) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_54_U43 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_54_n103), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_54_n133), .A(
        SD1_SB_inst_SD1_SB_bit_inst_54_n132), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_54_n134) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_54_U42 ( .A1(CipherErrorVec[94]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_54_n131), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_54_n130), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_54_n132) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_54_U41 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_54_n105), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_54_n99), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_54_n130) );
  OAI22_X1 SD1_SB_inst_SD1_SB_bit_inst_54_U40 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_54_n101), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_54_n129), .B1(CipherErrorVec[97]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_54_n128), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_54_n133) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_54_U39 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_54_n135), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_54_n136), .A(
        SD1_SB_inst_SD1_SB_bit_inst_54_n127), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_54_n138) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_54_U38 ( .A(StateRegOutput[54]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_54_n126), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_54_n127) );
  AOI211_X1 SD1_SB_inst_SD1_SB_bit_inst_54_U37 ( .C1(
        SD1_SB_inst_SD1_SB_bit_inst_54_n101), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_54_n125), .A(
        SD1_SB_inst_SD1_SB_bit_inst_54_n124), .B(
        SD1_SB_inst_SD1_SB_bit_inst_54_n123), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_54_n126) );
  AOI211_X1 SD1_SB_inst_SD1_SB_bit_inst_54_U36 ( .C1(
        SD1_SB_inst_SD1_SB_bit_inst_54_n122), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_54_n102), .A(
        SD1_SB_inst_SD1_SB_bit_inst_54_n121), .B(
        SD1_SB_inst_SD1_SB_bit_inst_54_n104), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_54_n123) );
  AOI22_X1 SD1_SB_inst_SD1_SB_bit_inst_54_U35 ( .A1(CipherErrorVec[91]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_54_n120), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_54_n99), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_54_n106), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_54_n122) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_54_U34 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_54_n102), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_54_n104), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_54_n119), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_54_n124) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_54_U33 ( .A(CipherErrorVec[97]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_54_n121) );
  OAI221_X1 SD1_SB_inst_SD1_SB_bit_inst_54_U32 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_54_n103), .B2(CipherErrorVec[97]), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_54_n103), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_54_n106), .A(CipherErrorVec[91]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_54_n118) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_54_U31 ( .A(StateRegOutput[52]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_54_n117), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_54_n136) );
  AOI22_X1 SD1_SB_inst_SD1_SB_bit_inst_54_U30 ( .A1(CipherErrorVec[94]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_54_n116), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_54_n101), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_54_n115), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_54_n117) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_54_U29 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_54_n103), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_54_n129), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_54_n115) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_54_U28 ( .A1(CipherErrorVec[91]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_54_n114), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_54_n129) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_54_U27 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_54_n120), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_54_n100), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_54_n114) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_54_U26 ( .A1(CipherErrorVec[94]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_54_n105), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_54_n120) );
  OAI21_X1 SD1_SB_inst_SD1_SB_bit_inst_54_U25 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_54_n131), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_54_n113), .A(
        SD1_SB_inst_SD1_SB_bit_inst_54_n128), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_54_n116) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_54_U24 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_54_n99), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_54_n106), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_54_n113) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_54_U23 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_54_n101), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_54_n103), .A3(CipherErrorVec[91]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_54_n131) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_54_U22 ( .A(StateRegOutput[55]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_54_n112), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_54_n135) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_54_U21 ( .B1(CipherErrorVec[97]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_54_n111), .A(
        SD1_SB_inst_SD1_SB_bit_inst_54_n110), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_54_n112) );
  AOI221_X1 SD1_SB_inst_SD1_SB_bit_inst_54_U20 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_54_n104), .B2(CipherErrorVec[91]), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_54_n102), .C2(CipherErrorVec[91]), .A(
        SD1_SB_inst_SD1_SB_bit_inst_54_n119), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_54_n110) );
  NAND3_X1 SD1_SB_inst_SD1_SB_bit_inst_54_U19 ( .A1(CipherErrorVec[94]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_54_n105), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_54_n99), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_54_n119) );
  OAI221_X1 SD1_SB_inst_SD1_SB_bit_inst_54_U18 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_54_n103), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_54_n128), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_54_n103), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_54_n109), .A(
        SD1_SB_inst_SD1_SB_bit_inst_54_n108), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_54_n111) );
  OAI21_X1 SD1_SB_inst_SD1_SB_bit_inst_54_U17 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_54_n105), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_54_n107), .A(CipherErrorVec[94]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_54_n108) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_54_U16 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_54_n101), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_54_n99), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_54_n104), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_54_n107) );
  OAI211_X1 SD1_SB_inst_SD1_SB_bit_inst_54_U15 ( .C1(CipherErrorVec[94]), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_54_n105), .A(
        SD1_SB_inst_SD1_SB_bit_inst_54_n99), .B(
        SD1_SB_inst_SD1_SB_bit_inst_54_n102), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_54_n109) );
  NAND3_X1 SD1_SB_inst_SD1_SB_bit_inst_54_U14 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_54_n101), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_54_n105), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_54_n100), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_54_n128) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_54_U13 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_54_n106), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_54_n105) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_54_U12 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_54_n104), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_54_n103) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_54_U11 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_54_n102), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_54_n101) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_54_U10 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_54_n100), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_54_n99) );
  MUX2_X1 SD1_SB_inst_SD1_SB_bit_inst_54_U9 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_54_n97), .B(
        SD1_SB_inst_SD1_SB_bit_inst_54_n98), .S(
        SD1_SB_inst_SD1_SB_bit_inst_54_n99), .Z(
        SD1_SB_inst_SD1_SB_bit_inst_54_n125) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_54_U8 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_54_n118), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_54_n97) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_54_U7 ( .A(CipherErrorVec[95]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_54_n104) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_54_U6 ( .A(CipherErrorVec[93]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_54_n102) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_54_U5 ( .A(CipherErrorVec[96]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_54_n106) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_54_U4 ( .A(CipherErrorVec[92]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_54_n100) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_54_U3 ( .A1(CipherErrorVec[94]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_54_n121), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_54_n98) );
  AOI222_X1 SD1_SB_inst_SD1_SB_bit_inst_55_U45 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_55_n141), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_55_n140), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_55_n141), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_55_n139), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_55_n140), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_55_n138), .ZN(Feedback[11]) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_55_U44 ( .A(StateRegOutput[52]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_55_n137), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_55_n138) );
  AOI211_X1 SD1_SB_inst_SD1_SB_bit_inst_55_U43 ( .C1(
        SD1_SB_inst_SD1_SB_bit_inst_55_n136), .C2(CipherErrorVec[94]), .A(
        SD1_SB_inst_SD1_SB_bit_inst_55_n135), .B(
        SD1_SB_inst_SD1_SB_bit_inst_55_n134), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_55_n137) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_55_U42 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_55_n105), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_55_n103), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_55_n133), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_55_n134) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_55_U41 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_55_n107), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_55_n132), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_55_n131), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_55_n135) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_55_U40 ( .A1(CipherErrorVec[94]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_55_n100), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_55_n131) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_55_U39 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_55_n130), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_55_n136) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_55_U38 ( .A(StateRegOutput[54]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_55_n129), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_55_n139) );
  AOI22_X1 SD1_SB_inst_SD1_SB_bit_inst_55_U37 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_55_n128), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_55_n127), .B1(CipherErrorVec[97]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_55_n126), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_55_n129) );
  OAI211_X1 SD1_SB_inst_SD1_SB_bit_inst_55_U36 ( .C1(
        SD1_SB_inst_SD1_SB_bit_inst_55_n125), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_55_n101), .A(
        SD1_SB_inst_SD1_SB_bit_inst_55_n124), .B(
        SD1_SB_inst_SD1_SB_bit_inst_55_n123), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_55_n126) );
  NAND3_X1 SD1_SB_inst_SD1_SB_bit_inst_55_U35 ( .A1(CipherErrorVec[91]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_55_n108), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_55_n122), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_55_n123) );
  OAI22_X1 SD1_SB_inst_SD1_SB_bit_inst_55_U34 ( .A1(CipherErrorVec[94]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_55_n106), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_55_n100), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_55_n103), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_55_n122) );
  AOI22_X1 SD1_SB_inst_SD1_SB_bit_inst_55_U33 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_55_n102), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_55_n104), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_55_n105), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_55_n108), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_55_n125) );
  OAI21_X1 SD1_SB_inst_SD1_SB_bit_inst_55_U32 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_55_n100), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_55_n121), .A(
        SD1_SB_inst_SD1_SB_bit_inst_55_n120), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_55_n127) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_55_U31 ( .A(CipherErrorVec[91]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_55_n121) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_55_U30 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_55_n124), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_55_n128) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_55_U29 ( .A(StateRegOutput[53]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_55_n119), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_55_n140) );
  AOI22_X1 SD1_SB_inst_SD1_SB_bit_inst_55_U28 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_55_n105), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_55_n118), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_55_n100), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_55_n117), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_55_n119) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_55_U27 ( .A1(CipherErrorVec[94]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_55_n132), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_55_n108), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_55_n117) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_55_U26 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_55_n102), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_55_n105), .A3(CipherErrorVec[91]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_55_n132) );
  OAI22_X1 SD1_SB_inst_SD1_SB_bit_inst_55_U25 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_55_n102), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_55_n133), .B1(CipherErrorVec[97]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_55_n130), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_55_n118) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_55_U24 ( .A1(CipherErrorVec[91]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_55_n116), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_55_n133) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_55_U23 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_55_n115), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_55_n101), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_55_n116) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_55_U22 ( .A1(CipherErrorVec[94]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_55_n107), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_55_n115) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_55_U21 ( .A(StateRegOutput[55]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_55_n114), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_55_n141) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_55_U20 ( .B1(CipherErrorVec[97]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_55_n113), .A(
        SD1_SB_inst_SD1_SB_bit_inst_55_n112), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_55_n114) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_55_U19 ( .B1(CipherErrorVec[91]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_55_n124), .A(
        SD1_SB_inst_SD1_SB_bit_inst_55_n120), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_55_n112) );
  NAND3_X1 SD1_SB_inst_SD1_SB_bit_inst_55_U18 ( .A1(CipherErrorVec[94]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_55_n100), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_55_n107), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_55_n120) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_55_U17 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_55_n102), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_55_n105), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_55_n124) );
  OAI221_X1 SD1_SB_inst_SD1_SB_bit_inst_55_U16 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_55_n105), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_55_n130), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_55_n105), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_55_n111), .A(
        SD1_SB_inst_SD1_SB_bit_inst_55_n110), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_55_n113) );
  OAI21_X1 SD1_SB_inst_SD1_SB_bit_inst_55_U15 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_55_n107), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_55_n109), .A(CipherErrorVec[94]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_55_n110) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_55_U14 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_55_n102), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_55_n100), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_55_n106), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_55_n109) );
  OAI211_X1 SD1_SB_inst_SD1_SB_bit_inst_55_U13 ( .C1(CipherErrorVec[94]), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_55_n107), .A(
        SD1_SB_inst_SD1_SB_bit_inst_55_n100), .B(
        SD1_SB_inst_SD1_SB_bit_inst_55_n103), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_55_n111) );
  NAND3_X1 SD1_SB_inst_SD1_SB_bit_inst_55_U12 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_55_n102), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_55_n107), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_55_n101), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_55_n130) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_55_U11 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_55_n108), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_55_n107) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_55_U10 ( .A(CipherErrorVec[95]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_55_n106) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_55_U9 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_55_n106), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_55_n105) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_55_U8 ( .A(CipherErrorVec[94]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_55_n104) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_55_U7 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_55_n103), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_55_n102) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_55_U6 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_55_n101), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_55_n100) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_55_U5 ( .A(CipherErrorVec[93]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_55_n103) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_55_U4 ( .A(CipherErrorVec[96]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_55_n108) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_55_U3 ( .A(CipherErrorVec[92]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_55_n101) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_56_U47 ( .B1(OutputRegIn[58]), .B2(
        OutputRegIn[59]), .A(SD1_SB_inst_SD1_SB_bit_inst_56_n131), .ZN(
        Feedback[12]) );
  AOI221_X1 SD1_SB_inst_SD1_SB_bit_inst_56_U46 ( .B1(OutputRegIn[58]), .B2(
        OutputRegIn[56]), .C1(OutputRegIn[59]), .C2(OutputRegIn[56]), .A(
        OutputRegIn[57]), .ZN(SD1_SB_inst_SD1_SB_bit_inst_56_n131) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_56_U45 ( .A(StateRegOutput[59]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_56_n127), .ZN(OutputRegIn[59]) );
  AOI211_X1 SD1_SB_inst_SD1_SB_bit_inst_56_U44 ( .C1(CipherErrorVec[104]), 
        .C2(SD1_SB_inst_SD1_SB_bit_inst_56_n126), .A(
        SD1_SB_inst_SD1_SB_bit_inst_56_n125), .B(
        SD1_SB_inst_SD1_SB_bit_inst_56_n124), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_56_n127) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_56_U43 ( .A1(CipherErrorVec[98]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_56_n101), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_56_n123), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_56_n124) );
  AOI222_X1 SD1_SB_inst_SD1_SB_bit_inst_56_U42 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_56_n108), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_56_n104), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_56_n108), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_56_n122), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_56_n104), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_56_n121), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_56_n126) );
  OAI221_X1 SD1_SB_inst_SD1_SB_bit_inst_56_U41 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_56_n120), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_56_n100), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_56_n120), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_56_n102), .A(
        SD1_SB_inst_SD1_SB_bit_inst_56_n106), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_56_n121) );
  OAI211_X1 SD1_SB_inst_SD1_SB_bit_inst_56_U40 ( .C1(
        SD1_SB_inst_SD1_SB_bit_inst_56_n105), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_56_n100), .A(
        SD1_SB_inst_SD1_SB_bit_inst_56_n119), .B(
        SD1_SB_inst_SD1_SB_bit_inst_56_n102), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_56_n122) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_56_U39 ( .A(StateRegOutput[58]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_56_n118), .ZN(OutputRegIn[58]) );
  AOI211_X1 SD1_SB_inst_SD1_SB_bit_inst_56_U38 ( .C1(CipherErrorVec[104]), 
        .C2(SD1_SB_inst_SD1_SB_bit_inst_56_n117), .A(
        SD1_SB_inst_SD1_SB_bit_inst_56_n125), .B(
        SD1_SB_inst_SD1_SB_bit_inst_56_n116), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_56_n118) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_56_U37 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_56_n128), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_56_n96), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_56_n116) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_56_U36 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_56_n105), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_56_n120), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_56_n128) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_56_U35 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_56_n102), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_56_n123), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_56_n119), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_56_n125) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_56_U34 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_56_n105), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_56_n100), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_56_n119) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_56_U33 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_56_n107), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_56_n103), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_56_n123) );
  OAI22_X1 SD1_SB_inst_SD1_SB_bit_inst_56_U32 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_56_n107), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_56_n115), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_56_n114), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_56_n102), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_56_n117) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_56_U31 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_56_n100), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_56_n104), .A(
        SD1_SB_inst_SD1_SB_bit_inst_56_n105), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_56_n114) );
  AOI22_X1 SD1_SB_inst_SD1_SB_bit_inst_56_U30 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_56_n105), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_56_n100), .B1(CipherErrorVec[98]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_56_n113), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_56_n115) );
  OAI21_X1 SD1_SB_inst_SD1_SB_bit_inst_56_U29 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_56_n103), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_56_n106), .A(
        SD1_SB_inst_SD1_SB_bit_inst_56_n112), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_56_n113) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_56_U28 ( .A(StateRegOutput[56]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_56_n111), .ZN(OutputRegIn[56]) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_56_U27 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_56_n110), .B2(CipherErrorVec[100]), .A(
        SD1_SB_inst_SD1_SB_bit_inst_56_n109), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_56_n111) );
  AOI221_X1 SD1_SB_inst_SD1_SB_bit_inst_56_U26 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_56_n107), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_56_n112), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_56_n108), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_56_n129), .A(
        SD1_SB_inst_SD1_SB_bit_inst_56_n104), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_56_n109) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_56_U25 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_56_n120), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_56_n112) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_56_U24 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_56_n100), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_56_n102), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_56_n120) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_56_U23 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_56_n130), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_56_n105), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_56_n110) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_56_U22 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_56_n108), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_56_n107) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_56_U21 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_56_n106), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_56_n105) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_56_U20 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_56_n104), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_56_n103) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_56_U19 ( .A(CipherErrorVec[100]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_56_n102) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_56_U18 ( .A(CipherErrorVec[99]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_56_n101) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_56_U17 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_56_n101), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_56_n100) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_56_U16 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_56_n99), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_56_n130) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_56_U15 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_56_n97), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_56_n129) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_56_U14 ( .A(CipherErrorVec[98]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_56_n96) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_56_U13 ( .A(CipherErrorVec[103]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_56_n108) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_56_U12 ( .A(CipherErrorVec[102]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_56_n106) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_56_U11 ( .A(CipherErrorVec[101]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_56_n104) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_56_U10 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_56_n100), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_56_n107), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_56_n98) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_56_U9 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_56_n98), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_56_n104), .A(
        SD1_SB_inst_SD1_SB_bit_inst_56_n96), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_56_n99) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_56_U8 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_56_n105), .A2(CipherErrorVec[100]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_56_n95) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_56_U7 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_56_n95), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_56_n96), .A(
        SD1_SB_inst_SD1_SB_bit_inst_56_n101), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_56_n97) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_56_U6 ( .A(StateRegOutput[57]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_56_n94), .ZN(OutputRegIn[57]) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_56_U5 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_56_n107), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_56_n92), .A(
        SD1_SB_inst_SD1_SB_bit_inst_56_n93), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_56_n94) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_56_U4 ( .A1(CipherErrorVec[100]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_56_n130), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_56_n106), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_56_n93) );
  OAI22_X1 SD1_SB_inst_SD1_SB_bit_inst_56_U3 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_56_n103), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_56_n129), .B1(CipherErrorVec[104]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_56_n128), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_56_n92) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_57_U37 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_57_n110), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_57_n109), .A(
        SD1_SB_inst_SD1_SB_bit_inst_57_n108), .ZN(Feedback[13]) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_57_U36 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_57_n107), .B2(StateRegOutput[56]), .A(
        SD1_SB_inst_SD1_SB_bit_inst_57_n106), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_57_n108) );
  OAI22_X1 SD1_SB_inst_SD1_SB_bit_inst_57_U35 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_57_n109), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_57_n110), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_57_n107), .B2(StateRegOutput[56]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_57_n106) );
  AOI22_X1 SD1_SB_inst_SD1_SB_bit_inst_57_U34 ( .A1(CipherErrorVec[98]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_57_n105), .B1(CipherErrorVec[101]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_57_n104), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_57_n107) );
  OAI21_X1 SD1_SB_inst_SD1_SB_bit_inst_57_U33 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_57_n103), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_57_n102), .A(
        SD1_SB_inst_SD1_SB_bit_inst_57_n101), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_57_n104) );
  NAND3_X1 SD1_SB_inst_SD1_SB_bit_inst_57_U32 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_57_n79), .A2(CipherErrorVec[103]), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_57_n78), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_57_n101) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_57_U31 ( .A1(CipherErrorVec[98]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_57_n79), .A3(CipherErrorVec[102]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_57_n103) );
  AOI211_X1 SD1_SB_inst_SD1_SB_bit_inst_57_U30 ( .C1(
        SD1_SB_inst_SD1_SB_bit_inst_57_n100), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_57_n78), .A(CipherErrorVec[102]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_57_n80), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_57_n105) );
  XOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_57_U29 ( .A(StateRegOutput[58]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_57_n99), .Z(
        SD1_SB_inst_SD1_SB_bit_inst_57_n109) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_57_U28 ( .B1(CipherErrorVec[104]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_57_n98), .A(
        SD1_SB_inst_SD1_SB_bit_inst_57_n97), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_57_n99) );
  AOI221_X1 SD1_SB_inst_SD1_SB_bit_inst_57_U27 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_57_n77), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_57_n96), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_57_n78), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_57_n95), .A(
        SD1_SB_inst_SD1_SB_bit_inst_57_n94), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_57_n97) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_57_U26 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_57_n93), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_57_n94) );
  OAI22_X1 SD1_SB_inst_SD1_SB_bit_inst_57_U25 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_57_n92), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_57_n80), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_57_n91), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_57_n82), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_57_n98) );
  AOI211_X1 SD1_SB_inst_SD1_SB_bit_inst_57_U24 ( .C1(CipherErrorVec[98]), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_57_n100), .A(
        SD1_SB_inst_SD1_SB_bit_inst_57_n79), .B(
        SD1_SB_inst_SD1_SB_bit_inst_57_n90), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_57_n91) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_57_U23 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_57_n102), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_57_n90) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_57_U22 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_57_n77), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_57_n83), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_57_n102) );
  AOI22_X1 SD1_SB_inst_SD1_SB_bit_inst_57_U21 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_57_n77), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_57_n81), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_57_n89), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_57_n83), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_57_n92) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_57_U20 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_57_n77), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_57_n95), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_57_n89) );
  XOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_57_U19 ( .A(StateRegOutput[59]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_57_n88), .Z(
        SD1_SB_inst_SD1_SB_bit_inst_57_n110) );
  OAI21_X1 SD1_SB_inst_SD1_SB_bit_inst_57_U18 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_57_n87), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_57_n96), .A(
        SD1_SB_inst_SD1_SB_bit_inst_57_n86), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_57_n88) );
  OAI221_X1 SD1_SB_inst_SD1_SB_bit_inst_57_U17 ( .B1(CipherErrorVec[102]), 
        .B2(SD1_SB_inst_SD1_SB_bit_inst_57_n85), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_57_n82), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_57_n84), .A(CipherErrorVec[104]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_57_n86) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_57_U16 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_57_n77), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_57_n79), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_57_n81), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_57_n84) );
  OAI33_X1 SD1_SB_inst_SD1_SB_bit_inst_57_U15 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_57_n79), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_57_n100), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_57_n78), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_57_n80), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_57_n83), .B3(
        SD1_SB_inst_SD1_SB_bit_inst_57_n77), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_57_n85) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_57_U14 ( .A1(CipherErrorVec[101]), .A2(
        CipherErrorVec[103]), .ZN(SD1_SB_inst_SD1_SB_bit_inst_57_n100) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_57_U13 ( .A1(CipherErrorVec[101]), .A2(
        CipherErrorVec[103]), .ZN(SD1_SB_inst_SD1_SB_bit_inst_57_n96) );
  AOI221_X1 SD1_SB_inst_SD1_SB_bit_inst_57_U12 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_57_n93), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_57_n77), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_57_n95), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_57_n77), .A(CipherErrorVec[104]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_57_n87) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_57_U11 ( .A(CipherErrorVec[98]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_57_n95) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_57_U10 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_57_n80), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_57_n82), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_57_n93) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_57_U9 ( .A(CipherErrorVec[101]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_57_n81) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_57_U8 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_57_n80), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_57_n79) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_57_U7 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_57_n78), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_57_n77) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_57_U6 ( .A(CipherErrorVec[102]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_57_n82) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_57_U5 ( .A(CipherErrorVec[103]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_57_n83) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_57_U4 ( .A(CipherErrorVec[100]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_57_n80) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_57_U3 ( .A(CipherErrorVec[99]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_57_n78) );
  OAI22_X1 SD1_SB_inst_SD1_SB_bit_inst_58_U45 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_58_n138), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_58_n137), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_58_n136), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_58_n135), .ZN(Feedback[14]) );
  XOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_58_U44 ( .A(StateRegOutput[57]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_58_n134), .Z(
        SD1_SB_inst_SD1_SB_bit_inst_58_n137) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_58_U43 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_58_n103), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_58_n133), .A(
        SD1_SB_inst_SD1_SB_bit_inst_58_n132), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_58_n134) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_58_U42 ( .A1(CipherErrorVec[101]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_58_n131), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_58_n130), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_58_n132) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_58_U41 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_58_n105), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_58_n99), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_58_n130) );
  OAI22_X1 SD1_SB_inst_SD1_SB_bit_inst_58_U40 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_58_n101), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_58_n129), .B1(CipherErrorVec[104]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_58_n128), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_58_n133) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_58_U39 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_58_n135), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_58_n136), .A(
        SD1_SB_inst_SD1_SB_bit_inst_58_n127), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_58_n138) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_58_U38 ( .A(StateRegOutput[58]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_58_n126), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_58_n127) );
  AOI211_X1 SD1_SB_inst_SD1_SB_bit_inst_58_U37 ( .C1(
        SD1_SB_inst_SD1_SB_bit_inst_58_n101), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_58_n125), .A(
        SD1_SB_inst_SD1_SB_bit_inst_58_n124), .B(
        SD1_SB_inst_SD1_SB_bit_inst_58_n123), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_58_n126) );
  AOI211_X1 SD1_SB_inst_SD1_SB_bit_inst_58_U36 ( .C1(
        SD1_SB_inst_SD1_SB_bit_inst_58_n122), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_58_n102), .A(
        SD1_SB_inst_SD1_SB_bit_inst_58_n121), .B(
        SD1_SB_inst_SD1_SB_bit_inst_58_n104), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_58_n123) );
  AOI22_X1 SD1_SB_inst_SD1_SB_bit_inst_58_U35 ( .A1(CipherErrorVec[98]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_58_n120), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_58_n99), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_58_n106), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_58_n122) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_58_U34 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_58_n102), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_58_n104), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_58_n119), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_58_n124) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_58_U33 ( .A(CipherErrorVec[104]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_58_n121) );
  OAI221_X1 SD1_SB_inst_SD1_SB_bit_inst_58_U32 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_58_n103), .B2(CipherErrorVec[104]), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_58_n103), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_58_n106), .A(CipherErrorVec[98]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_58_n118) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_58_U31 ( .A(StateRegOutput[56]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_58_n117), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_58_n136) );
  AOI22_X1 SD1_SB_inst_SD1_SB_bit_inst_58_U30 ( .A1(CipherErrorVec[101]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_58_n116), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_58_n101), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_58_n115), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_58_n117) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_58_U29 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_58_n103), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_58_n129), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_58_n115) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_58_U28 ( .A1(CipherErrorVec[98]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_58_n114), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_58_n129) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_58_U27 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_58_n120), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_58_n100), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_58_n114) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_58_U26 ( .A1(CipherErrorVec[101]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_58_n105), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_58_n120) );
  OAI21_X1 SD1_SB_inst_SD1_SB_bit_inst_58_U25 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_58_n131), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_58_n113), .A(
        SD1_SB_inst_SD1_SB_bit_inst_58_n128), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_58_n116) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_58_U24 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_58_n99), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_58_n106), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_58_n113) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_58_U23 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_58_n101), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_58_n103), .A3(CipherErrorVec[98]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_58_n131) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_58_U22 ( .A(StateRegOutput[59]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_58_n112), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_58_n135) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_58_U21 ( .B1(CipherErrorVec[104]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_58_n111), .A(
        SD1_SB_inst_SD1_SB_bit_inst_58_n110), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_58_n112) );
  AOI221_X1 SD1_SB_inst_SD1_SB_bit_inst_58_U20 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_58_n104), .B2(CipherErrorVec[98]), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_58_n102), .C2(CipherErrorVec[98]), .A(
        SD1_SB_inst_SD1_SB_bit_inst_58_n119), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_58_n110) );
  NAND3_X1 SD1_SB_inst_SD1_SB_bit_inst_58_U19 ( .A1(CipherErrorVec[101]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_58_n105), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_58_n99), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_58_n119) );
  OAI221_X1 SD1_SB_inst_SD1_SB_bit_inst_58_U18 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_58_n103), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_58_n128), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_58_n103), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_58_n109), .A(
        SD1_SB_inst_SD1_SB_bit_inst_58_n108), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_58_n111) );
  OAI21_X1 SD1_SB_inst_SD1_SB_bit_inst_58_U17 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_58_n105), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_58_n107), .A(CipherErrorVec[101]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_58_n108) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_58_U16 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_58_n101), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_58_n99), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_58_n104), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_58_n107) );
  OAI211_X1 SD1_SB_inst_SD1_SB_bit_inst_58_U15 ( .C1(CipherErrorVec[101]), 
        .C2(SD1_SB_inst_SD1_SB_bit_inst_58_n105), .A(
        SD1_SB_inst_SD1_SB_bit_inst_58_n99), .B(
        SD1_SB_inst_SD1_SB_bit_inst_58_n102), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_58_n109) );
  NAND3_X1 SD1_SB_inst_SD1_SB_bit_inst_58_U14 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_58_n101), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_58_n105), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_58_n100), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_58_n128) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_58_U13 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_58_n106), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_58_n105) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_58_U12 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_58_n104), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_58_n103) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_58_U11 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_58_n102), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_58_n101) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_58_U10 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_58_n100), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_58_n99) );
  MUX2_X1 SD1_SB_inst_SD1_SB_bit_inst_58_U9 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_58_n97), .B(
        SD1_SB_inst_SD1_SB_bit_inst_58_n98), .S(
        SD1_SB_inst_SD1_SB_bit_inst_58_n99), .Z(
        SD1_SB_inst_SD1_SB_bit_inst_58_n125) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_58_U8 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_58_n118), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_58_n97) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_58_U7 ( .A(CipherErrorVec[102]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_58_n104) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_58_U6 ( .A(CipherErrorVec[100]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_58_n102) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_58_U5 ( .A(CipherErrorVec[103]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_58_n106) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_58_U4 ( .A(CipherErrorVec[99]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_58_n100) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_58_U3 ( .A1(CipherErrorVec[101]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_58_n121), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_58_n98) );
  AOI222_X1 SD1_SB_inst_SD1_SB_bit_inst_59_U45 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_59_n141), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_59_n140), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_59_n141), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_59_n139), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_59_n140), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_59_n138), .ZN(Feedback[15]) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_59_U44 ( .A(StateRegOutput[56]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_59_n137), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_59_n138) );
  AOI211_X1 SD1_SB_inst_SD1_SB_bit_inst_59_U43 ( .C1(
        SD1_SB_inst_SD1_SB_bit_inst_59_n136), .C2(CipherErrorVec[101]), .A(
        SD1_SB_inst_SD1_SB_bit_inst_59_n135), .B(
        SD1_SB_inst_SD1_SB_bit_inst_59_n134), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_59_n137) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_59_U42 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_59_n105), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_59_n103), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_59_n133), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_59_n134) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_59_U41 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_59_n107), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_59_n132), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_59_n131), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_59_n135) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_59_U40 ( .A1(CipherErrorVec[101]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_59_n100), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_59_n131) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_59_U39 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_59_n130), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_59_n136) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_59_U38 ( .A(StateRegOutput[58]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_59_n129), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_59_n139) );
  AOI22_X1 SD1_SB_inst_SD1_SB_bit_inst_59_U37 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_59_n128), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_59_n127), .B1(CipherErrorVec[104]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_59_n126), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_59_n129) );
  OAI211_X1 SD1_SB_inst_SD1_SB_bit_inst_59_U36 ( .C1(
        SD1_SB_inst_SD1_SB_bit_inst_59_n125), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_59_n101), .A(
        SD1_SB_inst_SD1_SB_bit_inst_59_n124), .B(
        SD1_SB_inst_SD1_SB_bit_inst_59_n123), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_59_n126) );
  NAND3_X1 SD1_SB_inst_SD1_SB_bit_inst_59_U35 ( .A1(CipherErrorVec[98]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_59_n108), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_59_n122), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_59_n123) );
  OAI22_X1 SD1_SB_inst_SD1_SB_bit_inst_59_U34 ( .A1(CipherErrorVec[101]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_59_n106), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_59_n100), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_59_n103), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_59_n122) );
  AOI22_X1 SD1_SB_inst_SD1_SB_bit_inst_59_U33 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_59_n102), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_59_n104), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_59_n105), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_59_n108), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_59_n125) );
  OAI21_X1 SD1_SB_inst_SD1_SB_bit_inst_59_U32 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_59_n100), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_59_n121), .A(
        SD1_SB_inst_SD1_SB_bit_inst_59_n120), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_59_n127) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_59_U31 ( .A(CipherErrorVec[98]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_59_n121) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_59_U30 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_59_n124), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_59_n128) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_59_U29 ( .A(StateRegOutput[57]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_59_n119), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_59_n140) );
  AOI22_X1 SD1_SB_inst_SD1_SB_bit_inst_59_U28 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_59_n105), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_59_n118), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_59_n100), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_59_n117), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_59_n119) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_59_U27 ( .A1(CipherErrorVec[101]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_59_n132), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_59_n108), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_59_n117) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_59_U26 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_59_n102), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_59_n105), .A3(CipherErrorVec[98]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_59_n132) );
  OAI22_X1 SD1_SB_inst_SD1_SB_bit_inst_59_U25 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_59_n102), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_59_n133), .B1(CipherErrorVec[104]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_59_n130), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_59_n118) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_59_U24 ( .A1(CipherErrorVec[98]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_59_n116), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_59_n133) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_59_U23 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_59_n115), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_59_n101), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_59_n116) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_59_U22 ( .A1(CipherErrorVec[101]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_59_n107), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_59_n115) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_59_U21 ( .A(StateRegOutput[59]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_59_n114), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_59_n141) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_59_U20 ( .B1(CipherErrorVec[104]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_59_n113), .A(
        SD1_SB_inst_SD1_SB_bit_inst_59_n112), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_59_n114) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_59_U19 ( .B1(CipherErrorVec[98]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_59_n124), .A(
        SD1_SB_inst_SD1_SB_bit_inst_59_n120), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_59_n112) );
  NAND3_X1 SD1_SB_inst_SD1_SB_bit_inst_59_U18 ( .A1(CipherErrorVec[101]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_59_n100), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_59_n107), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_59_n120) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_59_U17 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_59_n102), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_59_n105), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_59_n124) );
  OAI221_X1 SD1_SB_inst_SD1_SB_bit_inst_59_U16 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_59_n105), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_59_n130), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_59_n105), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_59_n111), .A(
        SD1_SB_inst_SD1_SB_bit_inst_59_n110), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_59_n113) );
  OAI21_X1 SD1_SB_inst_SD1_SB_bit_inst_59_U15 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_59_n107), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_59_n109), .A(CipherErrorVec[101]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_59_n110) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_59_U14 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_59_n102), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_59_n100), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_59_n106), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_59_n109) );
  OAI211_X1 SD1_SB_inst_SD1_SB_bit_inst_59_U13 ( .C1(CipherErrorVec[101]), 
        .C2(SD1_SB_inst_SD1_SB_bit_inst_59_n107), .A(
        SD1_SB_inst_SD1_SB_bit_inst_59_n100), .B(
        SD1_SB_inst_SD1_SB_bit_inst_59_n103), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_59_n111) );
  NAND3_X1 SD1_SB_inst_SD1_SB_bit_inst_59_U12 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_59_n102), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_59_n107), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_59_n101), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_59_n130) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_59_U11 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_59_n108), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_59_n107) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_59_U10 ( .A(CipherErrorVec[102]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_59_n106) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_59_U9 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_59_n106), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_59_n105) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_59_U8 ( .A(CipherErrorVec[101]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_59_n104) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_59_U7 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_59_n103), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_59_n102) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_59_U6 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_59_n101), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_59_n100) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_59_U5 ( .A(CipherErrorVec[100]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_59_n103) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_59_U4 ( .A(CipherErrorVec[103]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_59_n108) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_59_U3 ( .A(CipherErrorVec[99]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_59_n101) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_60_U47 ( .B1(OutputRegIn[62]), .B2(
        OutputRegIn[63]), .A(SD1_SB_inst_SD1_SB_bit_inst_60_n131), .ZN(
        Feedback[0]) );
  AOI221_X1 SD1_SB_inst_SD1_SB_bit_inst_60_U46 ( .B1(OutputRegIn[62]), .B2(
        OutputRegIn[60]), .C1(OutputRegIn[63]), .C2(OutputRegIn[60]), .A(
        OutputRegIn[61]), .ZN(SD1_SB_inst_SD1_SB_bit_inst_60_n131) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_60_U45 ( .A(StateRegOutput[63]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_60_n127), .ZN(OutputRegIn[63]) );
  AOI211_X1 SD1_SB_inst_SD1_SB_bit_inst_60_U44 ( .C1(CipherErrorVec[111]), 
        .C2(SD1_SB_inst_SD1_SB_bit_inst_60_n126), .A(
        SD1_SB_inst_SD1_SB_bit_inst_60_n125), .B(
        SD1_SB_inst_SD1_SB_bit_inst_60_n124), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_60_n127) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_60_U43 ( .A1(CipherErrorVec[105]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_60_n101), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_60_n123), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_60_n124) );
  AOI222_X1 SD1_SB_inst_SD1_SB_bit_inst_60_U42 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_60_n108), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_60_n104), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_60_n108), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_60_n122), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_60_n104), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_60_n121), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_60_n126) );
  OAI221_X1 SD1_SB_inst_SD1_SB_bit_inst_60_U41 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_60_n120), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_60_n100), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_60_n120), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_60_n102), .A(
        SD1_SB_inst_SD1_SB_bit_inst_60_n106), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_60_n121) );
  OAI211_X1 SD1_SB_inst_SD1_SB_bit_inst_60_U40 ( .C1(
        SD1_SB_inst_SD1_SB_bit_inst_60_n105), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_60_n100), .A(
        SD1_SB_inst_SD1_SB_bit_inst_60_n119), .B(
        SD1_SB_inst_SD1_SB_bit_inst_60_n102), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_60_n122) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_60_U39 ( .A(StateRegOutput[62]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_60_n118), .ZN(OutputRegIn[62]) );
  AOI211_X1 SD1_SB_inst_SD1_SB_bit_inst_60_U38 ( .C1(CipherErrorVec[111]), 
        .C2(SD1_SB_inst_SD1_SB_bit_inst_60_n117), .A(
        SD1_SB_inst_SD1_SB_bit_inst_60_n125), .B(
        SD1_SB_inst_SD1_SB_bit_inst_60_n116), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_60_n118) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_60_U37 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_60_n128), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_60_n96), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_60_n116) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_60_U36 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_60_n105), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_60_n120), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_60_n128) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_60_U35 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_60_n102), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_60_n123), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_60_n119), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_60_n125) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_60_U34 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_60_n105), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_60_n100), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_60_n119) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_60_U33 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_60_n107), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_60_n103), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_60_n123) );
  OAI22_X1 SD1_SB_inst_SD1_SB_bit_inst_60_U32 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_60_n107), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_60_n115), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_60_n114), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_60_n102), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_60_n117) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_60_U31 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_60_n100), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_60_n104), .A(
        SD1_SB_inst_SD1_SB_bit_inst_60_n105), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_60_n114) );
  AOI22_X1 SD1_SB_inst_SD1_SB_bit_inst_60_U30 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_60_n105), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_60_n100), .B1(CipherErrorVec[105]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_60_n113), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_60_n115) );
  OAI21_X1 SD1_SB_inst_SD1_SB_bit_inst_60_U29 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_60_n103), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_60_n106), .A(
        SD1_SB_inst_SD1_SB_bit_inst_60_n112), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_60_n113) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_60_U28 ( .A(StateRegOutput[60]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_60_n111), .ZN(OutputRegIn[60]) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_60_U27 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_60_n110), .B2(CipherErrorVec[107]), .A(
        SD1_SB_inst_SD1_SB_bit_inst_60_n109), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_60_n111) );
  AOI221_X1 SD1_SB_inst_SD1_SB_bit_inst_60_U26 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_60_n107), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_60_n112), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_60_n108), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_60_n129), .A(
        SD1_SB_inst_SD1_SB_bit_inst_60_n104), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_60_n109) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_60_U25 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_60_n120), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_60_n112) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_60_U24 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_60_n100), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_60_n102), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_60_n120) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_60_U23 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_60_n130), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_60_n105), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_60_n110) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_60_U22 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_60_n108), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_60_n107) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_60_U21 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_60_n106), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_60_n105) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_60_U20 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_60_n104), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_60_n103) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_60_U19 ( .A(CipherErrorVec[107]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_60_n102) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_60_U18 ( .A(CipherErrorVec[106]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_60_n101) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_60_U17 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_60_n101), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_60_n100) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_60_U16 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_60_n99), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_60_n130) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_60_U15 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_60_n97), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_60_n129) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_60_U14 ( .A(CipherErrorVec[105]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_60_n96) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_60_U13 ( .A(CipherErrorVec[110]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_60_n108) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_60_U12 ( .A(CipherErrorVec[109]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_60_n106) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_60_U11 ( .A(CipherErrorVec[108]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_60_n104) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_60_U10 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_60_n100), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_60_n107), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_60_n98) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_60_U9 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_60_n98), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_60_n104), .A(
        SD1_SB_inst_SD1_SB_bit_inst_60_n96), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_60_n99) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_60_U8 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_60_n105), .A2(CipherErrorVec[107]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_60_n95) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_60_U7 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_60_n95), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_60_n96), .A(
        SD1_SB_inst_SD1_SB_bit_inst_60_n101), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_60_n97) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_60_U6 ( .A(StateRegOutput[61]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_60_n94), .ZN(OutputRegIn[61]) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_60_U5 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_60_n107), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_60_n92), .A(
        SD1_SB_inst_SD1_SB_bit_inst_60_n93), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_60_n94) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_60_U4 ( .A1(CipherErrorVec[107]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_60_n130), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_60_n106), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_60_n93) );
  OAI22_X1 SD1_SB_inst_SD1_SB_bit_inst_60_U3 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_60_n103), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_60_n129), .B1(CipherErrorVec[111]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_60_n128), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_60_n92) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_61_U37 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_61_n110), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_61_n109), .A(
        SD1_SB_inst_SD1_SB_bit_inst_61_n108), .ZN(Feedback[1]) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_61_U36 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_61_n107), .B2(StateRegOutput[60]), .A(
        SD1_SB_inst_SD1_SB_bit_inst_61_n106), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_61_n108) );
  OAI22_X1 SD1_SB_inst_SD1_SB_bit_inst_61_U35 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_61_n109), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_61_n110), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_61_n107), .B2(StateRegOutput[60]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_61_n106) );
  AOI22_X1 SD1_SB_inst_SD1_SB_bit_inst_61_U34 ( .A1(CipherErrorVec[105]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_61_n105), .B1(CipherErrorVec[108]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_61_n104), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_61_n107) );
  OAI21_X1 SD1_SB_inst_SD1_SB_bit_inst_61_U33 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_61_n103), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_61_n102), .A(
        SD1_SB_inst_SD1_SB_bit_inst_61_n101), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_61_n104) );
  NAND3_X1 SD1_SB_inst_SD1_SB_bit_inst_61_U32 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_61_n79), .A2(CipherErrorVec[110]), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_61_n78), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_61_n101) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_61_U31 ( .A1(CipherErrorVec[105]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_61_n79), .A3(CipherErrorVec[109]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_61_n103) );
  AOI211_X1 SD1_SB_inst_SD1_SB_bit_inst_61_U30 ( .C1(
        SD1_SB_inst_SD1_SB_bit_inst_61_n100), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_61_n78), .A(CipherErrorVec[109]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_61_n80), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_61_n105) );
  XOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_61_U29 ( .A(StateRegOutput[62]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_61_n99), .Z(
        SD1_SB_inst_SD1_SB_bit_inst_61_n109) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_61_U28 ( .B1(CipherErrorVec[111]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_61_n98), .A(
        SD1_SB_inst_SD1_SB_bit_inst_61_n97), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_61_n99) );
  AOI221_X1 SD1_SB_inst_SD1_SB_bit_inst_61_U27 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_61_n77), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_61_n96), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_61_n78), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_61_n95), .A(
        SD1_SB_inst_SD1_SB_bit_inst_61_n94), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_61_n97) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_61_U26 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_61_n93), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_61_n94) );
  OAI22_X1 SD1_SB_inst_SD1_SB_bit_inst_61_U25 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_61_n92), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_61_n80), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_61_n91), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_61_n82), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_61_n98) );
  AOI211_X1 SD1_SB_inst_SD1_SB_bit_inst_61_U24 ( .C1(CipherErrorVec[105]), 
        .C2(SD1_SB_inst_SD1_SB_bit_inst_61_n100), .A(
        SD1_SB_inst_SD1_SB_bit_inst_61_n79), .B(
        SD1_SB_inst_SD1_SB_bit_inst_61_n90), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_61_n91) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_61_U23 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_61_n102), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_61_n90) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_61_U22 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_61_n77), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_61_n83), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_61_n102) );
  AOI22_X1 SD1_SB_inst_SD1_SB_bit_inst_61_U21 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_61_n77), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_61_n81), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_61_n89), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_61_n83), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_61_n92) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_61_U20 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_61_n77), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_61_n95), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_61_n89) );
  XOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_61_U19 ( .A(StateRegOutput[63]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_61_n88), .Z(
        SD1_SB_inst_SD1_SB_bit_inst_61_n110) );
  OAI21_X1 SD1_SB_inst_SD1_SB_bit_inst_61_U18 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_61_n87), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_61_n96), .A(
        SD1_SB_inst_SD1_SB_bit_inst_61_n86), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_61_n88) );
  OAI221_X1 SD1_SB_inst_SD1_SB_bit_inst_61_U17 ( .B1(CipherErrorVec[109]), 
        .B2(SD1_SB_inst_SD1_SB_bit_inst_61_n85), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_61_n82), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_61_n84), .A(CipherErrorVec[111]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_61_n86) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_61_U16 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_61_n77), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_61_n79), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_61_n81), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_61_n84) );
  OAI33_X1 SD1_SB_inst_SD1_SB_bit_inst_61_U15 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_61_n79), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_61_n100), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_61_n78), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_61_n80), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_61_n83), .B3(
        SD1_SB_inst_SD1_SB_bit_inst_61_n77), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_61_n85) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_61_U14 ( .A1(CipherErrorVec[108]), .A2(
        CipherErrorVec[110]), .ZN(SD1_SB_inst_SD1_SB_bit_inst_61_n100) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_61_U13 ( .A1(CipherErrorVec[108]), .A2(
        CipherErrorVec[110]), .ZN(SD1_SB_inst_SD1_SB_bit_inst_61_n96) );
  AOI221_X1 SD1_SB_inst_SD1_SB_bit_inst_61_U12 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_61_n93), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_61_n77), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_61_n95), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_61_n77), .A(CipherErrorVec[111]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_61_n87) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_61_U11 ( .A(CipherErrorVec[105]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_61_n95) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_61_U10 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_61_n80), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_61_n82), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_61_n93) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_61_U9 ( .A(CipherErrorVec[108]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_61_n81) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_61_U8 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_61_n80), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_61_n79) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_61_U7 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_61_n78), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_61_n77) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_61_U6 ( .A(CipherErrorVec[109]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_61_n82) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_61_U5 ( .A(CipherErrorVec[110]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_61_n83) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_61_U4 ( .A(CipherErrorVec[107]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_61_n80) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_61_U3 ( .A(CipherErrorVec[106]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_61_n78) );
  OAI22_X1 SD1_SB_inst_SD1_SB_bit_inst_62_U45 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_62_n138), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_62_n137), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_62_n136), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_62_n135), .ZN(Feedback[2]) );
  XOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_62_U44 ( .A(StateRegOutput[61]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_62_n134), .Z(
        SD1_SB_inst_SD1_SB_bit_inst_62_n137) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_62_U43 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_62_n103), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_62_n133), .A(
        SD1_SB_inst_SD1_SB_bit_inst_62_n132), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_62_n134) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_62_U42 ( .A1(CipherErrorVec[108]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_62_n131), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_62_n130), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_62_n132) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_62_U41 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_62_n105), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_62_n99), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_62_n130) );
  OAI22_X1 SD1_SB_inst_SD1_SB_bit_inst_62_U40 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_62_n101), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_62_n129), .B1(CipherErrorVec[111]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_62_n128), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_62_n133) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_62_U39 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_62_n135), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_62_n136), .A(
        SD1_SB_inst_SD1_SB_bit_inst_62_n127), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_62_n138) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_62_U38 ( .A(StateRegOutput[62]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_62_n126), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_62_n127) );
  AOI211_X1 SD1_SB_inst_SD1_SB_bit_inst_62_U37 ( .C1(
        SD1_SB_inst_SD1_SB_bit_inst_62_n101), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_62_n125), .A(
        SD1_SB_inst_SD1_SB_bit_inst_62_n124), .B(
        SD1_SB_inst_SD1_SB_bit_inst_62_n123), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_62_n126) );
  AOI211_X1 SD1_SB_inst_SD1_SB_bit_inst_62_U36 ( .C1(
        SD1_SB_inst_SD1_SB_bit_inst_62_n122), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_62_n102), .A(
        SD1_SB_inst_SD1_SB_bit_inst_62_n121), .B(
        SD1_SB_inst_SD1_SB_bit_inst_62_n104), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_62_n123) );
  AOI22_X1 SD1_SB_inst_SD1_SB_bit_inst_62_U35 ( .A1(CipherErrorVec[105]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_62_n120), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_62_n99), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_62_n106), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_62_n122) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_62_U34 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_62_n102), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_62_n104), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_62_n119), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_62_n124) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_62_U33 ( .A(CipherErrorVec[111]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_62_n121) );
  OAI221_X1 SD1_SB_inst_SD1_SB_bit_inst_62_U32 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_62_n103), .B2(CipherErrorVec[111]), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_62_n103), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_62_n106), .A(CipherErrorVec[105]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_62_n118) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_62_U31 ( .A(StateRegOutput[60]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_62_n117), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_62_n136) );
  AOI22_X1 SD1_SB_inst_SD1_SB_bit_inst_62_U30 ( .A1(CipherErrorVec[108]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_62_n116), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_62_n101), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_62_n115), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_62_n117) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_62_U29 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_62_n103), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_62_n129), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_62_n115) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_62_U28 ( .A1(CipherErrorVec[105]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_62_n114), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_62_n129) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_62_U27 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_62_n120), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_62_n100), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_62_n114) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_62_U26 ( .A1(CipherErrorVec[108]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_62_n105), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_62_n120) );
  OAI21_X1 SD1_SB_inst_SD1_SB_bit_inst_62_U25 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_62_n131), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_62_n113), .A(
        SD1_SB_inst_SD1_SB_bit_inst_62_n128), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_62_n116) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_62_U24 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_62_n99), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_62_n106), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_62_n113) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_62_U23 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_62_n101), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_62_n103), .A3(CipherErrorVec[105]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_62_n131) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_62_U22 ( .A(StateRegOutput[63]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_62_n112), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_62_n135) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_62_U21 ( .B1(CipherErrorVec[111]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_62_n111), .A(
        SD1_SB_inst_SD1_SB_bit_inst_62_n110), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_62_n112) );
  AOI221_X1 SD1_SB_inst_SD1_SB_bit_inst_62_U20 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_62_n104), .B2(CipherErrorVec[105]), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_62_n102), .C2(CipherErrorVec[105]), .A(
        SD1_SB_inst_SD1_SB_bit_inst_62_n119), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_62_n110) );
  NAND3_X1 SD1_SB_inst_SD1_SB_bit_inst_62_U19 ( .A1(CipherErrorVec[108]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_62_n105), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_62_n99), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_62_n119) );
  OAI221_X1 SD1_SB_inst_SD1_SB_bit_inst_62_U18 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_62_n103), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_62_n128), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_62_n103), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_62_n109), .A(
        SD1_SB_inst_SD1_SB_bit_inst_62_n108), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_62_n111) );
  OAI21_X1 SD1_SB_inst_SD1_SB_bit_inst_62_U17 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_62_n105), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_62_n107), .A(CipherErrorVec[108]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_62_n108) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_62_U16 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_62_n101), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_62_n99), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_62_n104), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_62_n107) );
  OAI211_X1 SD1_SB_inst_SD1_SB_bit_inst_62_U15 ( .C1(CipherErrorVec[108]), 
        .C2(SD1_SB_inst_SD1_SB_bit_inst_62_n105), .A(
        SD1_SB_inst_SD1_SB_bit_inst_62_n99), .B(
        SD1_SB_inst_SD1_SB_bit_inst_62_n102), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_62_n109) );
  NAND3_X1 SD1_SB_inst_SD1_SB_bit_inst_62_U14 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_62_n101), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_62_n105), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_62_n100), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_62_n128) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_62_U13 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_62_n106), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_62_n105) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_62_U12 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_62_n104), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_62_n103) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_62_U11 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_62_n102), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_62_n101) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_62_U10 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_62_n100), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_62_n99) );
  MUX2_X1 SD1_SB_inst_SD1_SB_bit_inst_62_U9 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_62_n97), .B(
        SD1_SB_inst_SD1_SB_bit_inst_62_n98), .S(
        SD1_SB_inst_SD1_SB_bit_inst_62_n99), .Z(
        SD1_SB_inst_SD1_SB_bit_inst_62_n125) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_62_U8 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_62_n118), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_62_n97) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_62_U7 ( .A(CipherErrorVec[109]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_62_n104) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_62_U6 ( .A(CipherErrorVec[107]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_62_n102) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_62_U5 ( .A(CipherErrorVec[110]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_62_n106) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_62_U4 ( .A(CipherErrorVec[106]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_62_n100) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_62_U3 ( .A1(CipherErrorVec[108]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_62_n121), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_62_n98) );
  AOI222_X1 SD1_SB_inst_SD1_SB_bit_inst_63_U45 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_63_n141), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_63_n140), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_63_n141), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_63_n139), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_63_n140), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_63_n138), .ZN(Feedback[3]) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_63_U44 ( .A(StateRegOutput[60]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_63_n137), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_63_n138) );
  AOI211_X1 SD1_SB_inst_SD1_SB_bit_inst_63_U43 ( .C1(
        SD1_SB_inst_SD1_SB_bit_inst_63_n136), .C2(CipherErrorVec[108]), .A(
        SD1_SB_inst_SD1_SB_bit_inst_63_n135), .B(
        SD1_SB_inst_SD1_SB_bit_inst_63_n134), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_63_n137) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_63_U42 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_63_n105), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_63_n103), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_63_n133), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_63_n134) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_63_U41 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_63_n107), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_63_n132), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_63_n131), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_63_n135) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_63_U40 ( .A1(CipherErrorVec[108]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_63_n100), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_63_n131) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_63_U39 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_63_n130), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_63_n136) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_63_U38 ( .A(StateRegOutput[62]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_63_n129), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_63_n139) );
  AOI22_X1 SD1_SB_inst_SD1_SB_bit_inst_63_U37 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_63_n128), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_63_n127), .B1(CipherErrorVec[111]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_63_n126), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_63_n129) );
  OAI211_X1 SD1_SB_inst_SD1_SB_bit_inst_63_U36 ( .C1(
        SD1_SB_inst_SD1_SB_bit_inst_63_n125), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_63_n101), .A(
        SD1_SB_inst_SD1_SB_bit_inst_63_n124), .B(
        SD1_SB_inst_SD1_SB_bit_inst_63_n123), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_63_n126) );
  NAND3_X1 SD1_SB_inst_SD1_SB_bit_inst_63_U35 ( .A1(CipherErrorVec[105]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_63_n108), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_63_n122), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_63_n123) );
  OAI22_X1 SD1_SB_inst_SD1_SB_bit_inst_63_U34 ( .A1(CipherErrorVec[108]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_63_n106), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_63_n100), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_63_n103), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_63_n122) );
  AOI22_X1 SD1_SB_inst_SD1_SB_bit_inst_63_U33 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_63_n102), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_63_n104), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_63_n105), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_63_n108), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_63_n125) );
  OAI21_X1 SD1_SB_inst_SD1_SB_bit_inst_63_U32 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_63_n100), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_63_n121), .A(
        SD1_SB_inst_SD1_SB_bit_inst_63_n120), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_63_n127) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_63_U31 ( .A(CipherErrorVec[105]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_63_n121) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_63_U30 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_63_n124), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_63_n128) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_63_U29 ( .A(StateRegOutput[61]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_63_n119), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_63_n140) );
  AOI22_X1 SD1_SB_inst_SD1_SB_bit_inst_63_U28 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_63_n105), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_63_n118), .B1(
        SD1_SB_inst_SD1_SB_bit_inst_63_n100), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_63_n117), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_63_n119) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_63_U27 ( .A1(CipherErrorVec[108]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_63_n132), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_63_n108), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_63_n117) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_63_U26 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_63_n102), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_63_n105), .A3(CipherErrorVec[105]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_63_n132) );
  OAI22_X1 SD1_SB_inst_SD1_SB_bit_inst_63_U25 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_63_n102), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_63_n133), .B1(CipherErrorVec[111]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_63_n130), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_63_n118) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_63_U24 ( .A1(CipherErrorVec[105]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_63_n116), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_63_n133) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_63_U23 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_63_n115), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_63_n101), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_63_n116) );
  NOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_63_U22 ( .A1(CipherErrorVec[108]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_63_n107), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_63_n115) );
  XNOR2_X1 SD1_SB_inst_SD1_SB_bit_inst_63_U21 ( .A(StateRegOutput[63]), .B(
        SD1_SB_inst_SD1_SB_bit_inst_63_n114), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_63_n141) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_63_U20 ( .B1(CipherErrorVec[111]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_63_n113), .A(
        SD1_SB_inst_SD1_SB_bit_inst_63_n112), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_63_n114) );
  AOI21_X1 SD1_SB_inst_SD1_SB_bit_inst_63_U19 ( .B1(CipherErrorVec[105]), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_63_n124), .A(
        SD1_SB_inst_SD1_SB_bit_inst_63_n120), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_63_n112) );
  NAND3_X1 SD1_SB_inst_SD1_SB_bit_inst_63_U18 ( .A1(CipherErrorVec[108]), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_63_n100), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_63_n107), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_63_n120) );
  NAND2_X1 SD1_SB_inst_SD1_SB_bit_inst_63_U17 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_63_n102), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_63_n105), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_63_n124) );
  OAI221_X1 SD1_SB_inst_SD1_SB_bit_inst_63_U16 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_63_n105), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_63_n130), .C1(
        SD1_SB_inst_SD1_SB_bit_inst_63_n105), .C2(
        SD1_SB_inst_SD1_SB_bit_inst_63_n111), .A(
        SD1_SB_inst_SD1_SB_bit_inst_63_n110), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_63_n113) );
  OAI21_X1 SD1_SB_inst_SD1_SB_bit_inst_63_U15 ( .B1(
        SD1_SB_inst_SD1_SB_bit_inst_63_n107), .B2(
        SD1_SB_inst_SD1_SB_bit_inst_63_n109), .A(CipherErrorVec[108]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_63_n110) );
  NOR3_X1 SD1_SB_inst_SD1_SB_bit_inst_63_U14 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_63_n102), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_63_n100), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_63_n106), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_63_n109) );
  OAI211_X1 SD1_SB_inst_SD1_SB_bit_inst_63_U13 ( .C1(CipherErrorVec[108]), 
        .C2(SD1_SB_inst_SD1_SB_bit_inst_63_n107), .A(
        SD1_SB_inst_SD1_SB_bit_inst_63_n100), .B(
        SD1_SB_inst_SD1_SB_bit_inst_63_n103), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_63_n111) );
  NAND3_X1 SD1_SB_inst_SD1_SB_bit_inst_63_U12 ( .A1(
        SD1_SB_inst_SD1_SB_bit_inst_63_n102), .A2(
        SD1_SB_inst_SD1_SB_bit_inst_63_n107), .A3(
        SD1_SB_inst_SD1_SB_bit_inst_63_n101), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_63_n130) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_63_U11 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_63_n108), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_63_n107) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_63_U10 ( .A(CipherErrorVec[109]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_63_n106) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_63_U9 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_63_n106), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_63_n105) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_63_U8 ( .A(CipherErrorVec[108]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_63_n104) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_63_U7 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_63_n103), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_63_n102) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_63_U6 ( .A(
        SD1_SB_inst_SD1_SB_bit_inst_63_n101), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_63_n100) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_63_U5 ( .A(CipherErrorVec[107]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_63_n103) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_63_U4 ( .A(CipherErrorVec[110]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_63_n108) );
  INV_X1 SD1_SB_inst_SD1_SB_bit_inst_63_U3 ( .A(CipherErrorVec[106]), .ZN(
        SD1_SB_inst_SD1_SB_bit_inst_63_n101) );
  XNOR2_X1 Red_PlaintextInst_LFInst_0_LFInst_0_U2 ( .A(
        Red_PlaintextInst_LFInst_0_LFInst_0_n3), .B(Input[2]), .ZN(
        Red_Input[0]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_0_LFInst_0_U1 ( .A(Input[0]), .B(Input[1]), 
        .ZN(Red_PlaintextInst_LFInst_0_LFInst_0_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_0_LFInst_1_U2 ( .A(
        Red_PlaintextInst_LFInst_0_LFInst_1_n3), .B(Input[3]), .ZN(
        Red_Input[1]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_0_LFInst_1_U1 ( .A(Input[0]), .B(Input[1]), 
        .ZN(Red_PlaintextInst_LFInst_0_LFInst_1_n3) );
  XOR2_X1 Red_PlaintextInst_LFInst_0_LFInst_2_U1 ( .A(Input[0]), .B(Input[2]), 
        .Z(Red_Input[2]) );
  XOR2_X1 Red_PlaintextInst_LFInst_0_LFInst_3_U1 ( .A(Input[0]), .B(Input[3]), 
        .Z(Red_Input[3]) );
  XOR2_X1 Red_PlaintextInst_LFInst_0_LFInst_4_U1 ( .A(Input[1]), .B(Input[2]), 
        .Z(Red_Input[4]) );
  XOR2_X1 Red_PlaintextInst_LFInst_0_LFInst_5_U1 ( .A(Input[1]), .B(Input[3]), 
        .Z(Red_Input[5]) );
  XOR2_X1 Red_PlaintextInst_LFInst_0_LFInst_6_U1 ( .A(Input[2]), .B(Input[3]), 
        .Z(Red_Input[6]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_1_LFInst_0_U2 ( .A(
        Red_PlaintextInst_LFInst_1_LFInst_0_n3), .B(Input[6]), .ZN(
        Red_Input[7]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_1_LFInst_0_U1 ( .A(Input[4]), .B(Input[5]), 
        .ZN(Red_PlaintextInst_LFInst_1_LFInst_0_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_1_LFInst_1_U2 ( .A(
        Red_PlaintextInst_LFInst_1_LFInst_1_n3), .B(Input[7]), .ZN(
        Red_Input[8]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_1_LFInst_1_U1 ( .A(Input[4]), .B(Input[5]), 
        .ZN(Red_PlaintextInst_LFInst_1_LFInst_1_n3) );
  XOR2_X1 Red_PlaintextInst_LFInst_1_LFInst_2_U1 ( .A(Input[4]), .B(Input[6]), 
        .Z(Red_Input[9]) );
  XOR2_X1 Red_PlaintextInst_LFInst_1_LFInst_3_U1 ( .A(Input[4]), .B(Input[7]), 
        .Z(Red_Input[10]) );
  XOR2_X1 Red_PlaintextInst_LFInst_1_LFInst_4_U1 ( .A(Input[5]), .B(Input[6]), 
        .Z(Red_Input[11]) );
  XOR2_X1 Red_PlaintextInst_LFInst_1_LFInst_5_U1 ( .A(Input[5]), .B(Input[7]), 
        .Z(Red_Input[12]) );
  XOR2_X1 Red_PlaintextInst_LFInst_1_LFInst_6_U1 ( .A(Input[6]), .B(Input[7]), 
        .Z(Red_Input[13]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_2_LFInst_0_U2 ( .A(
        Red_PlaintextInst_LFInst_2_LFInst_0_n3), .B(Input[10]), .ZN(
        Red_Input[14]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_2_LFInst_0_U1 ( .A(Input[8]), .B(Input[9]), 
        .ZN(Red_PlaintextInst_LFInst_2_LFInst_0_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_2_LFInst_1_U2 ( .A(
        Red_PlaintextInst_LFInst_2_LFInst_1_n3), .B(Input[11]), .ZN(
        Red_Input[15]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_2_LFInst_1_U1 ( .A(Input[8]), .B(Input[9]), 
        .ZN(Red_PlaintextInst_LFInst_2_LFInst_1_n3) );
  XOR2_X1 Red_PlaintextInst_LFInst_2_LFInst_2_U1 ( .A(Input[8]), .B(Input[10]), 
        .Z(Red_Input[16]) );
  XOR2_X1 Red_PlaintextInst_LFInst_2_LFInst_3_U1 ( .A(Input[8]), .B(Input[11]), 
        .Z(Red_Input[17]) );
  XOR2_X1 Red_PlaintextInst_LFInst_2_LFInst_4_U1 ( .A(Input[9]), .B(Input[10]), 
        .Z(Red_Input[18]) );
  XOR2_X1 Red_PlaintextInst_LFInst_2_LFInst_5_U1 ( .A(Input[9]), .B(Input[11]), 
        .Z(Red_Input[19]) );
  XOR2_X1 Red_PlaintextInst_LFInst_2_LFInst_6_U1 ( .A(Input[10]), .B(Input[11]), .Z(Red_Input[20]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_3_LFInst_0_U2 ( .A(
        Red_PlaintextInst_LFInst_3_LFInst_0_n3), .B(Input[14]), .ZN(
        Red_Input[21]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_3_LFInst_0_U1 ( .A(Input[12]), .B(
        Input[13]), .ZN(Red_PlaintextInst_LFInst_3_LFInst_0_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_3_LFInst_1_U2 ( .A(
        Red_PlaintextInst_LFInst_3_LFInst_1_n3), .B(Input[15]), .ZN(
        Red_Input[22]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_3_LFInst_1_U1 ( .A(Input[12]), .B(
        Input[13]), .ZN(Red_PlaintextInst_LFInst_3_LFInst_1_n3) );
  XOR2_X1 Red_PlaintextInst_LFInst_3_LFInst_2_U1 ( .A(Input[12]), .B(Input[14]), .Z(Red_Input[23]) );
  XOR2_X1 Red_PlaintextInst_LFInst_3_LFInst_3_U1 ( .A(Input[12]), .B(Input[15]), .Z(Red_Input[24]) );
  XOR2_X1 Red_PlaintextInst_LFInst_3_LFInst_4_U1 ( .A(Input[13]), .B(Input[14]), .Z(Red_Input[25]) );
  XOR2_X1 Red_PlaintextInst_LFInst_3_LFInst_5_U1 ( .A(Input[13]), .B(Input[15]), .Z(Red_Input[26]) );
  XOR2_X1 Red_PlaintextInst_LFInst_3_LFInst_6_U1 ( .A(Input[14]), .B(Input[15]), .Z(Red_Input[27]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_4_LFInst_0_U2 ( .A(
        Red_PlaintextInst_LFInst_4_LFInst_0_n3), .B(Input[18]), .ZN(
        Red_Input[28]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_4_LFInst_0_U1 ( .A(Input[16]), .B(
        Input[17]), .ZN(Red_PlaintextInst_LFInst_4_LFInst_0_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_4_LFInst_1_U2 ( .A(
        Red_PlaintextInst_LFInst_4_LFInst_1_n3), .B(Input[19]), .ZN(
        Red_Input[29]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_4_LFInst_1_U1 ( .A(Input[16]), .B(
        Input[17]), .ZN(Red_PlaintextInst_LFInst_4_LFInst_1_n3) );
  XOR2_X1 Red_PlaintextInst_LFInst_4_LFInst_2_U1 ( .A(Input[16]), .B(Input[18]), .Z(Red_Input[30]) );
  XOR2_X1 Red_PlaintextInst_LFInst_4_LFInst_3_U1 ( .A(Input[16]), .B(Input[19]), .Z(Red_Input[31]) );
  XOR2_X1 Red_PlaintextInst_LFInst_4_LFInst_4_U1 ( .A(Input[17]), .B(Input[18]), .Z(Red_Input[32]) );
  XOR2_X1 Red_PlaintextInst_LFInst_4_LFInst_5_U1 ( .A(Input[17]), .B(Input[19]), .Z(Red_Input[33]) );
  XOR2_X1 Red_PlaintextInst_LFInst_4_LFInst_6_U1 ( .A(Input[18]), .B(Input[19]), .Z(Red_Input[34]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_5_LFInst_0_U2 ( .A(
        Red_PlaintextInst_LFInst_5_LFInst_0_n3), .B(Input[22]), .ZN(
        Red_Input[35]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_5_LFInst_0_U1 ( .A(Input[20]), .B(
        Input[21]), .ZN(Red_PlaintextInst_LFInst_5_LFInst_0_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_5_LFInst_1_U2 ( .A(
        Red_PlaintextInst_LFInst_5_LFInst_1_n3), .B(Input[23]), .ZN(
        Red_Input[36]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_5_LFInst_1_U1 ( .A(Input[20]), .B(
        Input[21]), .ZN(Red_PlaintextInst_LFInst_5_LFInst_1_n3) );
  XOR2_X1 Red_PlaintextInst_LFInst_5_LFInst_2_U1 ( .A(Input[20]), .B(Input[22]), .Z(Red_Input[37]) );
  XOR2_X1 Red_PlaintextInst_LFInst_5_LFInst_3_U1 ( .A(Input[20]), .B(Input[23]), .Z(Red_Input[38]) );
  XOR2_X1 Red_PlaintextInst_LFInst_5_LFInst_4_U1 ( .A(Input[21]), .B(Input[22]), .Z(Red_Input[39]) );
  XOR2_X1 Red_PlaintextInst_LFInst_5_LFInst_5_U1 ( .A(Input[21]), .B(Input[23]), .Z(Red_Input[40]) );
  XOR2_X1 Red_PlaintextInst_LFInst_5_LFInst_6_U1 ( .A(Input[22]), .B(Input[23]), .Z(Red_Input[41]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_6_LFInst_0_U2 ( .A(
        Red_PlaintextInst_LFInst_6_LFInst_0_n3), .B(Input[26]), .ZN(
        Red_Input[42]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_6_LFInst_0_U1 ( .A(Input[24]), .B(
        Input[25]), .ZN(Red_PlaintextInst_LFInst_6_LFInst_0_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_6_LFInst_1_U2 ( .A(
        Red_PlaintextInst_LFInst_6_LFInst_1_n3), .B(Input[27]), .ZN(
        Red_Input[43]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_6_LFInst_1_U1 ( .A(Input[24]), .B(
        Input[25]), .ZN(Red_PlaintextInst_LFInst_6_LFInst_1_n3) );
  XOR2_X1 Red_PlaintextInst_LFInst_6_LFInst_2_U1 ( .A(Input[24]), .B(Input[26]), .Z(Red_Input[44]) );
  XOR2_X1 Red_PlaintextInst_LFInst_6_LFInst_3_U1 ( .A(Input[24]), .B(Input[27]), .Z(Red_Input[45]) );
  XOR2_X1 Red_PlaintextInst_LFInst_6_LFInst_4_U1 ( .A(Input[25]), .B(Input[26]), .Z(Red_Input[46]) );
  XOR2_X1 Red_PlaintextInst_LFInst_6_LFInst_5_U1 ( .A(Input[25]), .B(Input[27]), .Z(Red_Input[47]) );
  XOR2_X1 Red_PlaintextInst_LFInst_6_LFInst_6_U1 ( .A(Input[26]), .B(Input[27]), .Z(Red_Input[48]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_7_LFInst_0_U2 ( .A(
        Red_PlaintextInst_LFInst_7_LFInst_0_n3), .B(Input[30]), .ZN(
        Red_Input[49]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_7_LFInst_0_U1 ( .A(Input[28]), .B(
        Input[29]), .ZN(Red_PlaintextInst_LFInst_7_LFInst_0_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_7_LFInst_1_U2 ( .A(
        Red_PlaintextInst_LFInst_7_LFInst_1_n3), .B(Input[31]), .ZN(
        Red_Input[50]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_7_LFInst_1_U1 ( .A(Input[28]), .B(
        Input[29]), .ZN(Red_PlaintextInst_LFInst_7_LFInst_1_n3) );
  XOR2_X1 Red_PlaintextInst_LFInst_7_LFInst_2_U1 ( .A(Input[28]), .B(Input[30]), .Z(Red_Input[51]) );
  XOR2_X1 Red_PlaintextInst_LFInst_7_LFInst_3_U1 ( .A(Input[28]), .B(Input[31]), .Z(Red_Input[52]) );
  XOR2_X1 Red_PlaintextInst_LFInst_7_LFInst_4_U1 ( .A(Input[29]), .B(Input[30]), .Z(Red_Input[53]) );
  XOR2_X1 Red_PlaintextInst_LFInst_7_LFInst_5_U1 ( .A(Input[29]), .B(Input[31]), .Z(Red_Input[54]) );
  XOR2_X1 Red_PlaintextInst_LFInst_7_LFInst_6_U1 ( .A(Input[30]), .B(Input[31]), .Z(Red_Input[55]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_8_LFInst_0_U2 ( .A(
        Red_PlaintextInst_LFInst_8_LFInst_0_n3), .B(Input[34]), .ZN(
        Red_Input[56]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_8_LFInst_0_U1 ( .A(Input[32]), .B(
        Input[33]), .ZN(Red_PlaintextInst_LFInst_8_LFInst_0_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_8_LFInst_1_U2 ( .A(
        Red_PlaintextInst_LFInst_8_LFInst_1_n3), .B(Input[35]), .ZN(
        Red_Input[57]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_8_LFInst_1_U1 ( .A(Input[32]), .B(
        Input[33]), .ZN(Red_PlaintextInst_LFInst_8_LFInst_1_n3) );
  XOR2_X1 Red_PlaintextInst_LFInst_8_LFInst_2_U1 ( .A(Input[32]), .B(Input[34]), .Z(Red_Input[58]) );
  XOR2_X1 Red_PlaintextInst_LFInst_8_LFInst_3_U1 ( .A(Input[32]), .B(Input[35]), .Z(Red_Input[59]) );
  XOR2_X1 Red_PlaintextInst_LFInst_8_LFInst_4_U1 ( .A(Input[33]), .B(Input[34]), .Z(Red_Input[60]) );
  XOR2_X1 Red_PlaintextInst_LFInst_8_LFInst_5_U1 ( .A(Input[33]), .B(Input[35]), .Z(Red_Input[61]) );
  XOR2_X1 Red_PlaintextInst_LFInst_8_LFInst_6_U1 ( .A(Input[34]), .B(Input[35]), .Z(Red_Input[62]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_9_LFInst_0_U2 ( .A(
        Red_PlaintextInst_LFInst_9_LFInst_0_n3), .B(Input[38]), .ZN(
        Red_Input[63]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_9_LFInst_0_U1 ( .A(Input[36]), .B(
        Input[37]), .ZN(Red_PlaintextInst_LFInst_9_LFInst_0_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_9_LFInst_1_U2 ( .A(
        Red_PlaintextInst_LFInst_9_LFInst_1_n3), .B(Input[39]), .ZN(
        Red_Input[64]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_9_LFInst_1_U1 ( .A(Input[36]), .B(
        Input[37]), .ZN(Red_PlaintextInst_LFInst_9_LFInst_1_n3) );
  XOR2_X1 Red_PlaintextInst_LFInst_9_LFInst_2_U1 ( .A(Input[36]), .B(Input[38]), .Z(Red_Input[65]) );
  XOR2_X1 Red_PlaintextInst_LFInst_9_LFInst_3_U1 ( .A(Input[36]), .B(Input[39]), .Z(Red_Input[66]) );
  XOR2_X1 Red_PlaintextInst_LFInst_9_LFInst_4_U1 ( .A(Input[37]), .B(Input[38]), .Z(Red_Input[67]) );
  XOR2_X1 Red_PlaintextInst_LFInst_9_LFInst_5_U1 ( .A(Input[37]), .B(Input[39]), .Z(Red_Input[68]) );
  XOR2_X1 Red_PlaintextInst_LFInst_9_LFInst_6_U1 ( .A(Input[38]), .B(Input[39]), .Z(Red_Input[69]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_10_LFInst_0_U2 ( .A(
        Red_PlaintextInst_LFInst_10_LFInst_0_n3), .B(Input[42]), .ZN(
        Red_Input[70]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_10_LFInst_0_U1 ( .A(Input[40]), .B(
        Input[41]), .ZN(Red_PlaintextInst_LFInst_10_LFInst_0_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_10_LFInst_1_U2 ( .A(
        Red_PlaintextInst_LFInst_10_LFInst_1_n3), .B(Input[43]), .ZN(
        Red_Input[71]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_10_LFInst_1_U1 ( .A(Input[40]), .B(
        Input[41]), .ZN(Red_PlaintextInst_LFInst_10_LFInst_1_n3) );
  XOR2_X1 Red_PlaintextInst_LFInst_10_LFInst_2_U1 ( .A(Input[40]), .B(
        Input[42]), .Z(Red_Input[72]) );
  XOR2_X1 Red_PlaintextInst_LFInst_10_LFInst_3_U1 ( .A(Input[40]), .B(
        Input[43]), .Z(Red_Input[73]) );
  XOR2_X1 Red_PlaintextInst_LFInst_10_LFInst_4_U1 ( .A(Input[41]), .B(
        Input[42]), .Z(Red_Input[74]) );
  XOR2_X1 Red_PlaintextInst_LFInst_10_LFInst_5_U1 ( .A(Input[41]), .B(
        Input[43]), .Z(Red_Input[75]) );
  XOR2_X1 Red_PlaintextInst_LFInst_10_LFInst_6_U1 ( .A(Input[42]), .B(
        Input[43]), .Z(Red_Input[76]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_11_LFInst_0_U2 ( .A(
        Red_PlaintextInst_LFInst_11_LFInst_0_n3), .B(Input[46]), .ZN(
        Red_Input[77]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_11_LFInst_0_U1 ( .A(Input[44]), .B(
        Input[45]), .ZN(Red_PlaintextInst_LFInst_11_LFInst_0_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_11_LFInst_1_U2 ( .A(
        Red_PlaintextInst_LFInst_11_LFInst_1_n3), .B(Input[47]), .ZN(
        Red_Input[78]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_11_LFInst_1_U1 ( .A(Input[44]), .B(
        Input[45]), .ZN(Red_PlaintextInst_LFInst_11_LFInst_1_n3) );
  XOR2_X1 Red_PlaintextInst_LFInst_11_LFInst_2_U1 ( .A(Input[44]), .B(
        Input[46]), .Z(Red_Input[79]) );
  XOR2_X1 Red_PlaintextInst_LFInst_11_LFInst_3_U1 ( .A(Input[44]), .B(
        Input[47]), .Z(Red_Input[80]) );
  XOR2_X1 Red_PlaintextInst_LFInst_11_LFInst_4_U1 ( .A(Input[45]), .B(
        Input[46]), .Z(Red_Input[81]) );
  XOR2_X1 Red_PlaintextInst_LFInst_11_LFInst_5_U1 ( .A(Input[45]), .B(
        Input[47]), .Z(Red_Input[82]) );
  XOR2_X1 Red_PlaintextInst_LFInst_11_LFInst_6_U1 ( .A(Input[46]), .B(
        Input[47]), .Z(Red_Input[83]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_12_LFInst_0_U2 ( .A(
        Red_PlaintextInst_LFInst_12_LFInst_0_n3), .B(Input[50]), .ZN(
        Red_Input[84]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_12_LFInst_0_U1 ( .A(Input[48]), .B(
        Input[49]), .ZN(Red_PlaintextInst_LFInst_12_LFInst_0_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_12_LFInst_1_U2 ( .A(
        Red_PlaintextInst_LFInst_12_LFInst_1_n3), .B(Input[51]), .ZN(
        Red_Input[85]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_12_LFInst_1_U1 ( .A(Input[48]), .B(
        Input[49]), .ZN(Red_PlaintextInst_LFInst_12_LFInst_1_n3) );
  XOR2_X1 Red_PlaintextInst_LFInst_12_LFInst_2_U1 ( .A(Input[48]), .B(
        Input[50]), .Z(Red_Input[86]) );
  XOR2_X1 Red_PlaintextInst_LFInst_12_LFInst_3_U1 ( .A(Input[48]), .B(
        Input[51]), .Z(Red_Input[87]) );
  XOR2_X1 Red_PlaintextInst_LFInst_12_LFInst_4_U1 ( .A(Input[49]), .B(
        Input[50]), .Z(Red_Input[88]) );
  XOR2_X1 Red_PlaintextInst_LFInst_12_LFInst_5_U1 ( .A(Input[49]), .B(
        Input[51]), .Z(Red_Input[89]) );
  XOR2_X1 Red_PlaintextInst_LFInst_12_LFInst_6_U1 ( .A(Input[50]), .B(
        Input[51]), .Z(Red_Input[90]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_13_LFInst_0_U2 ( .A(
        Red_PlaintextInst_LFInst_13_LFInst_0_n3), .B(Input[54]), .ZN(
        Red_Input[91]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_13_LFInst_0_U1 ( .A(Input[52]), .B(
        Input[53]), .ZN(Red_PlaintextInst_LFInst_13_LFInst_0_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_13_LFInst_1_U2 ( .A(
        Red_PlaintextInst_LFInst_13_LFInst_1_n3), .B(Input[55]), .ZN(
        Red_Input[92]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_13_LFInst_1_U1 ( .A(Input[52]), .B(
        Input[53]), .ZN(Red_PlaintextInst_LFInst_13_LFInst_1_n3) );
  XOR2_X1 Red_PlaintextInst_LFInst_13_LFInst_2_U1 ( .A(Input[52]), .B(
        Input[54]), .Z(Red_Input[93]) );
  XOR2_X1 Red_PlaintextInst_LFInst_13_LFInst_3_U1 ( .A(Input[52]), .B(
        Input[55]), .Z(Red_Input[94]) );
  XOR2_X1 Red_PlaintextInst_LFInst_13_LFInst_4_U1 ( .A(Input[53]), .B(
        Input[54]), .Z(Red_Input[95]) );
  XOR2_X1 Red_PlaintextInst_LFInst_13_LFInst_5_U1 ( .A(Input[53]), .B(
        Input[55]), .Z(Red_Input[96]) );
  XOR2_X1 Red_PlaintextInst_LFInst_13_LFInst_6_U1 ( .A(Input[54]), .B(
        Input[55]), .Z(Red_Input[97]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_14_LFInst_0_U2 ( .A(
        Red_PlaintextInst_LFInst_14_LFInst_0_n3), .B(Input[58]), .ZN(
        Red_Input[98]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_14_LFInst_0_U1 ( .A(Input[56]), .B(
        Input[57]), .ZN(Red_PlaintextInst_LFInst_14_LFInst_0_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_14_LFInst_1_U2 ( .A(
        Red_PlaintextInst_LFInst_14_LFInst_1_n3), .B(Input[59]), .ZN(
        Red_Input[99]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_14_LFInst_1_U1 ( .A(Input[56]), .B(
        Input[57]), .ZN(Red_PlaintextInst_LFInst_14_LFInst_1_n3) );
  XOR2_X1 Red_PlaintextInst_LFInst_14_LFInst_2_U1 ( .A(Input[56]), .B(
        Input[58]), .Z(Red_Input[100]) );
  XOR2_X1 Red_PlaintextInst_LFInst_14_LFInst_3_U1 ( .A(Input[56]), .B(
        Input[59]), .Z(Red_Input[101]) );
  XOR2_X1 Red_PlaintextInst_LFInst_14_LFInst_4_U1 ( .A(Input[57]), .B(
        Input[58]), .Z(Red_Input[102]) );
  XOR2_X1 Red_PlaintextInst_LFInst_14_LFInst_5_U1 ( .A(Input[57]), .B(
        Input[59]), .Z(Red_Input[103]) );
  XOR2_X1 Red_PlaintextInst_LFInst_14_LFInst_6_U1 ( .A(Input[58]), .B(
        Input[59]), .Z(Red_Input[104]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_15_LFInst_0_U2 ( .A(
        Red_PlaintextInst_LFInst_15_LFInst_0_n3), .B(Input[62]), .ZN(
        Red_Input[105]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_15_LFInst_0_U1 ( .A(Input[60]), .B(
        Input[61]), .ZN(Red_PlaintextInst_LFInst_15_LFInst_0_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_15_LFInst_1_U2 ( .A(
        Red_PlaintextInst_LFInst_15_LFInst_1_n3), .B(Input[63]), .ZN(
        Red_Input[106]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_15_LFInst_1_U1 ( .A(Input[60]), .B(
        Input[61]), .ZN(Red_PlaintextInst_LFInst_15_LFInst_1_n3) );
  XOR2_X1 Red_PlaintextInst_LFInst_15_LFInst_2_U1 ( .A(Input[60]), .B(
        Input[62]), .Z(Red_Input[107]) );
  XOR2_X1 Red_PlaintextInst_LFInst_15_LFInst_3_U1 ( .A(Input[60]), .B(
        Input[63]), .Z(Red_Input[108]) );
  XOR2_X1 Red_PlaintextInst_LFInst_15_LFInst_4_U1 ( .A(Input[61]), .B(
        Input[62]), .Z(Red_Input[109]) );
  XOR2_X1 Red_PlaintextInst_LFInst_15_LFInst_5_U1 ( .A(Input[61]), .B(
        Input[63]), .Z(Red_Input[110]) );
  XOR2_X1 Red_PlaintextInst_LFInst_15_LFInst_6_U1 ( .A(Input[62]), .B(
        Input[63]), .Z(Red_Input[111]) );
  MUX2_X1 Red_InputMUX_MUXInst_0_U1 ( .A(Red_Feedback[0]), .B(Red_Input[0]), 
        .S(rst), .Z(Red_MCOutput[0]) );
  MUX2_X1 Red_InputMUX_MUXInst_1_U1 ( .A(Red_Feedback[1]), .B(Red_Input[1]), 
        .S(rst), .Z(Red_MCOutput[1]) );
  MUX2_X1 Red_InputMUX_MUXInst_2_U1 ( .A(Red_Feedback[2]), .B(Red_Input[2]), 
        .S(rst), .Z(Red_MCOutput[2]) );
  MUX2_X1 Red_InputMUX_MUXInst_3_U1 ( .A(Red_Feedback[3]), .B(Red_Input[3]), 
        .S(rst), .Z(Red_MCOutput[3]) );
  MUX2_X1 Red_InputMUX_MUXInst_4_U1 ( .A(Red_Feedback[4]), .B(Red_Input[4]), 
        .S(rst), .Z(Red_MCOutput[4]) );
  MUX2_X1 Red_InputMUX_MUXInst_5_U1 ( .A(Red_Feedback[5]), .B(Red_Input[5]), 
        .S(rst), .Z(Red_MCOutput[5]) );
  MUX2_X1 Red_InputMUX_MUXInst_6_U1 ( .A(Red_Feedback[6]), .B(Red_Input[6]), 
        .S(rst), .Z(Red_MCOutput[6]) );
  MUX2_X1 Red_InputMUX_MUXInst_7_U1 ( .A(Red_Feedback[7]), .B(Red_Input[7]), 
        .S(rst), .Z(Red_MCOutput[7]) );
  MUX2_X1 Red_InputMUX_MUXInst_8_U1 ( .A(Red_Feedback[8]), .B(Red_Input[8]), 
        .S(rst), .Z(Red_MCOutput[8]) );
  MUX2_X1 Red_InputMUX_MUXInst_9_U1 ( .A(Red_Feedback[9]), .B(Red_Input[9]), 
        .S(rst), .Z(Red_MCOutput[9]) );
  MUX2_X1 Red_InputMUX_MUXInst_10_U1 ( .A(Red_Feedback[10]), .B(Red_Input[10]), 
        .S(rst), .Z(Red_MCOutput[10]) );
  MUX2_X1 Red_InputMUX_MUXInst_11_U1 ( .A(Red_Feedback[11]), .B(Red_Input[11]), 
        .S(rst), .Z(Red_MCOutput[11]) );
  MUX2_X1 Red_InputMUX_MUXInst_12_U1 ( .A(Red_Feedback[12]), .B(Red_Input[12]), 
        .S(rst), .Z(Red_MCOutput[12]) );
  MUX2_X1 Red_InputMUX_MUXInst_13_U1 ( .A(Red_Feedback[13]), .B(Red_Input[13]), 
        .S(rst), .Z(Red_MCOutput[13]) );
  MUX2_X1 Red_InputMUX_MUXInst_14_U1 ( .A(Red_Feedback[14]), .B(Red_Input[14]), 
        .S(rst), .Z(Red_MCOutput[14]) );
  MUX2_X1 Red_InputMUX_MUXInst_15_U1 ( .A(Red_Feedback[15]), .B(Red_Input[15]), 
        .S(rst), .Z(Red_MCOutput[15]) );
  MUX2_X1 Red_InputMUX_MUXInst_16_U1 ( .A(Red_Feedback[16]), .B(Red_Input[16]), 
        .S(rst), .Z(Red_MCOutput[16]) );
  MUX2_X1 Red_InputMUX_MUXInst_17_U1 ( .A(Red_Feedback[17]), .B(Red_Input[17]), 
        .S(rst), .Z(Red_MCOutput[17]) );
  MUX2_X1 Red_InputMUX_MUXInst_18_U1 ( .A(Red_Feedback[18]), .B(Red_Input[18]), 
        .S(rst), .Z(Red_MCOutput[18]) );
  MUX2_X1 Red_InputMUX_MUXInst_19_U1 ( .A(Red_Feedback[19]), .B(Red_Input[19]), 
        .S(rst), .Z(Red_MCOutput[19]) );
  MUX2_X1 Red_InputMUX_MUXInst_20_U1 ( .A(Red_Feedback[20]), .B(Red_Input[20]), 
        .S(rst), .Z(Red_MCOutput[20]) );
  MUX2_X1 Red_InputMUX_MUXInst_21_U1 ( .A(Red_Feedback[21]), .B(Red_Input[21]), 
        .S(rst), .Z(Red_MCOutput[21]) );
  MUX2_X1 Red_InputMUX_MUXInst_22_U1 ( .A(Red_Feedback[22]), .B(Red_Input[22]), 
        .S(rst), .Z(Red_MCOutput[22]) );
  MUX2_X1 Red_InputMUX_MUXInst_23_U1 ( .A(Red_Feedback[23]), .B(Red_Input[23]), 
        .S(rst), .Z(Red_MCOutput[23]) );
  MUX2_X1 Red_InputMUX_MUXInst_24_U1 ( .A(Red_Feedback[24]), .B(Red_Input[24]), 
        .S(rst), .Z(Red_MCOutput[24]) );
  MUX2_X1 Red_InputMUX_MUXInst_25_U1 ( .A(Red_Feedback[25]), .B(Red_Input[25]), 
        .S(rst), .Z(Red_MCOutput[25]) );
  MUX2_X1 Red_InputMUX_MUXInst_26_U1 ( .A(Red_Feedback[26]), .B(Red_Input[26]), 
        .S(rst), .Z(Red_MCOutput[26]) );
  MUX2_X1 Red_InputMUX_MUXInst_27_U1 ( .A(Red_Feedback[27]), .B(Red_Input[27]), 
        .S(rst), .Z(Red_MCOutput[27]) );
  MUX2_X1 Red_InputMUX_MUXInst_28_U1 ( .A(Red_Feedback[28]), .B(Red_Input[28]), 
        .S(rst), .Z(Red_MCOutput[28]) );
  MUX2_X1 Red_InputMUX_MUXInst_29_U1 ( .A(Red_Feedback[29]), .B(Red_Input[29]), 
        .S(rst), .Z(Red_MCOutput[29]) );
  MUX2_X1 Red_InputMUX_MUXInst_30_U1 ( .A(Red_Feedback[30]), .B(Red_Input[30]), 
        .S(rst), .Z(Red_MCOutput[30]) );
  MUX2_X1 Red_InputMUX_MUXInst_31_U1 ( .A(Red_Feedback[31]), .B(Red_Input[31]), 
        .S(rst), .Z(Red_MCOutput[31]) );
  MUX2_X1 Red_InputMUX_MUXInst_32_U1 ( .A(Red_Feedback[32]), .B(Red_Input[32]), 
        .S(rst), .Z(Red_MCOutput[32]) );
  MUX2_X1 Red_InputMUX_MUXInst_33_U1 ( .A(Red_Feedback[33]), .B(Red_Input[33]), 
        .S(rst), .Z(Red_MCOutput[33]) );
  MUX2_X1 Red_InputMUX_MUXInst_34_U1 ( .A(Red_Feedback[34]), .B(Red_Input[34]), 
        .S(rst), .Z(Red_MCOutput[34]) );
  MUX2_X1 Red_InputMUX_MUXInst_35_U1 ( .A(Red_Feedback[35]), .B(Red_Input[35]), 
        .S(rst), .Z(Red_MCOutput[35]) );
  MUX2_X1 Red_InputMUX_MUXInst_36_U1 ( .A(Red_Feedback[36]), .B(Red_Input[36]), 
        .S(rst), .Z(Red_MCOutput[36]) );
  MUX2_X1 Red_InputMUX_MUXInst_37_U1 ( .A(Red_Feedback[37]), .B(Red_Input[37]), 
        .S(rst), .Z(Red_MCOutput[37]) );
  MUX2_X1 Red_InputMUX_MUXInst_38_U1 ( .A(Red_Feedback[38]), .B(Red_Input[38]), 
        .S(rst), .Z(Red_MCOutput[38]) );
  MUX2_X1 Red_InputMUX_MUXInst_39_U1 ( .A(Red_Feedback[39]), .B(Red_Input[39]), 
        .S(rst), .Z(Red_MCOutput[39]) );
  MUX2_X1 Red_InputMUX_MUXInst_40_U1 ( .A(Red_Feedback[40]), .B(Red_Input[40]), 
        .S(rst), .Z(Red_MCOutput[40]) );
  MUX2_X1 Red_InputMUX_MUXInst_41_U1 ( .A(Red_Feedback[41]), .B(Red_Input[41]), 
        .S(rst), .Z(Red_MCOutput[41]) );
  MUX2_X1 Red_InputMUX_MUXInst_42_U1 ( .A(Red_Feedback[42]), .B(Red_Input[42]), 
        .S(rst), .Z(Red_MCOutput[42]) );
  MUX2_X1 Red_InputMUX_MUXInst_43_U1 ( .A(Red_Feedback[43]), .B(Red_Input[43]), 
        .S(rst), .Z(Red_MCOutput[43]) );
  MUX2_X1 Red_InputMUX_MUXInst_44_U1 ( .A(Red_Feedback[44]), .B(Red_Input[44]), 
        .S(rst), .Z(Red_MCOutput[44]) );
  MUX2_X1 Red_InputMUX_MUXInst_45_U1 ( .A(Red_Feedback[45]), .B(Red_Input[45]), 
        .S(rst), .Z(Red_MCOutput[45]) );
  MUX2_X1 Red_InputMUX_MUXInst_46_U1 ( .A(Red_Feedback[46]), .B(Red_Input[46]), 
        .S(rst), .Z(Red_MCOutput[46]) );
  MUX2_X1 Red_InputMUX_MUXInst_47_U1 ( .A(Red_Feedback[47]), .B(Red_Input[47]), 
        .S(rst), .Z(Red_MCOutput[47]) );
  MUX2_X1 Red_InputMUX_MUXInst_48_U1 ( .A(Red_Feedback[48]), .B(Red_Input[48]), 
        .S(rst), .Z(Red_MCOutput[48]) );
  MUX2_X1 Red_InputMUX_MUXInst_49_U1 ( .A(Red_Feedback[49]), .B(Red_Input[49]), 
        .S(rst), .Z(Red_MCOutput[49]) );
  MUX2_X1 Red_InputMUX_MUXInst_50_U1 ( .A(Red_Feedback[50]), .B(Red_Input[50]), 
        .S(rst), .Z(Red_MCOutput[50]) );
  MUX2_X1 Red_InputMUX_MUXInst_51_U1 ( .A(Red_Feedback[51]), .B(Red_Input[51]), 
        .S(rst), .Z(Red_MCOutput[51]) );
  MUX2_X1 Red_InputMUX_MUXInst_52_U1 ( .A(Red_Feedback[52]), .B(Red_Input[52]), 
        .S(rst), .Z(Red_MCOutput[52]) );
  MUX2_X1 Red_InputMUX_MUXInst_53_U1 ( .A(Red_Feedback[53]), .B(Red_Input[53]), 
        .S(rst), .Z(Red_MCOutput[53]) );
  MUX2_X1 Red_InputMUX_MUXInst_54_U1 ( .A(Red_Feedback[54]), .B(Red_Input[54]), 
        .S(rst), .Z(Red_MCOutput[54]) );
  MUX2_X1 Red_InputMUX_MUXInst_55_U1 ( .A(Red_Feedback[55]), .B(Red_Input[55]), 
        .S(rst), .Z(Red_MCOutput[55]) );
  MUX2_X1 Red_InputMUX_MUXInst_56_U1 ( .A(Red_Feedback[56]), .B(Red_Input[56]), 
        .S(rst), .Z(Red_MCInput[56]) );
  MUX2_X1 Red_InputMUX_MUXInst_57_U1 ( .A(Red_Feedback[57]), .B(Red_Input[57]), 
        .S(rst), .Z(Red_MCInput[57]) );
  MUX2_X1 Red_InputMUX_MUXInst_58_U1 ( .A(Red_Feedback[58]), .B(Red_Input[58]), 
        .S(rst), .Z(Red_MCInput[58]) );
  MUX2_X1 Red_InputMUX_MUXInst_59_U1 ( .A(Red_Feedback[59]), .B(Red_Input[59]), 
        .S(rst), .Z(Red_MCInput[59]) );
  MUX2_X1 Red_InputMUX_MUXInst_60_U1 ( .A(Red_Feedback[60]), .B(Red_Input[60]), 
        .S(rst), .Z(Red_MCInput[60]) );
  MUX2_X1 Red_InputMUX_MUXInst_61_U1 ( .A(Red_Feedback[61]), .B(Red_Input[61]), 
        .S(rst), .Z(Red_MCInput[61]) );
  MUX2_X1 Red_InputMUX_MUXInst_62_U1 ( .A(Red_Feedback[62]), .B(Red_Input[62]), 
        .S(rst), .Z(Red_MCInput[62]) );
  MUX2_X1 Red_InputMUX_MUXInst_63_U1 ( .A(Red_Feedback[63]), .B(Red_Input[63]), 
        .S(rst), .Z(Red_MCInput[63]) );
  MUX2_X1 Red_InputMUX_MUXInst_64_U1 ( .A(Red_Feedback[64]), .B(Red_Input[64]), 
        .S(rst), .Z(Red_MCInput[64]) );
  MUX2_X1 Red_InputMUX_MUXInst_65_U1 ( .A(Red_Feedback[65]), .B(Red_Input[65]), 
        .S(rst), .Z(Red_MCInput[65]) );
  MUX2_X1 Red_InputMUX_MUXInst_66_U1 ( .A(Red_Feedback[66]), .B(Red_Input[66]), 
        .S(rst), .Z(Red_MCInput[66]) );
  MUX2_X1 Red_InputMUX_MUXInst_67_U1 ( .A(Red_Feedback[67]), .B(Red_Input[67]), 
        .S(rst), .Z(Red_MCInput[67]) );
  MUX2_X1 Red_InputMUX_MUXInst_68_U1 ( .A(Red_Feedback[68]), .B(Red_Input[68]), 
        .S(rst), .Z(Red_MCInput[68]) );
  MUX2_X1 Red_InputMUX_MUXInst_69_U1 ( .A(Red_Feedback[69]), .B(Red_Input[69]), 
        .S(rst), .Z(Red_MCInput[69]) );
  MUX2_X1 Red_InputMUX_MUXInst_70_U1 ( .A(Red_Feedback[70]), .B(Red_Input[70]), 
        .S(rst), .Z(Red_MCInput[70]) );
  MUX2_X1 Red_InputMUX_MUXInst_71_U1 ( .A(Red_Feedback[71]), .B(Red_Input[71]), 
        .S(rst), .Z(Red_MCInput[71]) );
  MUX2_X1 Red_InputMUX_MUXInst_72_U1 ( .A(Red_Feedback[72]), .B(Red_Input[72]), 
        .S(rst), .Z(Red_MCInput[72]) );
  MUX2_X1 Red_InputMUX_MUXInst_73_U1 ( .A(Red_Feedback[73]), .B(Red_Input[73]), 
        .S(rst), .Z(Red_MCInput[73]) );
  MUX2_X1 Red_InputMUX_MUXInst_74_U1 ( .A(Red_Feedback[74]), .B(Red_Input[74]), 
        .S(rst), .Z(Red_MCInput[74]) );
  MUX2_X1 Red_InputMUX_MUXInst_75_U1 ( .A(Red_Feedback[75]), .B(Red_Input[75]), 
        .S(rst), .Z(Red_MCInput[75]) );
  MUX2_X1 Red_InputMUX_MUXInst_76_U1 ( .A(Red_Feedback[76]), .B(Red_Input[76]), 
        .S(rst), .Z(Red_MCInput[76]) );
  MUX2_X1 Red_InputMUX_MUXInst_77_U1 ( .A(Red_Feedback[77]), .B(Red_Input[77]), 
        .S(rst), .Z(Red_MCInput[77]) );
  MUX2_X1 Red_InputMUX_MUXInst_78_U1 ( .A(Red_Feedback[78]), .B(Red_Input[78]), 
        .S(rst), .Z(Red_MCInput[78]) );
  MUX2_X1 Red_InputMUX_MUXInst_79_U1 ( .A(Red_Feedback[79]), .B(Red_Input[79]), 
        .S(rst), .Z(Red_MCInput[79]) );
  MUX2_X1 Red_InputMUX_MUXInst_80_U1 ( .A(Red_Feedback[80]), .B(Red_Input[80]), 
        .S(rst), .Z(Red_MCInput[80]) );
  MUX2_X1 Red_InputMUX_MUXInst_81_U1 ( .A(Red_Feedback[81]), .B(Red_Input[81]), 
        .S(rst), .Z(Red_MCInput[81]) );
  MUX2_X1 Red_InputMUX_MUXInst_82_U1 ( .A(Red_Feedback[82]), .B(Red_Input[82]), 
        .S(rst), .Z(Red_MCInput[82]) );
  MUX2_X1 Red_InputMUX_MUXInst_83_U1 ( .A(Red_Feedback[83]), .B(Red_Input[83]), 
        .S(rst), .Z(Red_MCInput[83]) );
  MUX2_X1 Red_InputMUX_MUXInst_84_U1 ( .A(Red_Feedback[84]), .B(Red_Input[84]), 
        .S(rst), .Z(Red_MCInput[84]) );
  MUX2_X1 Red_InputMUX_MUXInst_85_U1 ( .A(Red_Feedback[85]), .B(Red_Input[85]), 
        .S(rst), .Z(Red_MCInput[85]) );
  MUX2_X1 Red_InputMUX_MUXInst_86_U1 ( .A(Red_Feedback[86]), .B(Red_Input[86]), 
        .S(rst), .Z(Red_MCInput[86]) );
  MUX2_X1 Red_InputMUX_MUXInst_87_U1 ( .A(Red_Feedback[87]), .B(Red_Input[87]), 
        .S(rst), .Z(Red_MCInput[87]) );
  MUX2_X1 Red_InputMUX_MUXInst_88_U1 ( .A(Red_Feedback[88]), .B(Red_Input[88]), 
        .S(rst), .Z(Red_MCInput[88]) );
  MUX2_X1 Red_InputMUX_MUXInst_89_U1 ( .A(Red_Feedback[89]), .B(Red_Input[89]), 
        .S(rst), .Z(Red_MCInput[89]) );
  MUX2_X1 Red_InputMUX_MUXInst_90_U1 ( .A(Red_Feedback[90]), .B(Red_Input[90]), 
        .S(rst), .Z(Red_MCInput[90]) );
  MUX2_X1 Red_InputMUX_MUXInst_91_U1 ( .A(Red_Feedback[91]), .B(Red_Input[91]), 
        .S(rst), .Z(Red_MCInput[91]) );
  MUX2_X1 Red_InputMUX_MUXInst_92_U1 ( .A(Red_Feedback[92]), .B(Red_Input[92]), 
        .S(rst), .Z(Red_MCInput[92]) );
  MUX2_X1 Red_InputMUX_MUXInst_93_U1 ( .A(Red_Feedback[93]), .B(Red_Input[93]), 
        .S(rst), .Z(Red_MCInput[93]) );
  MUX2_X1 Red_InputMUX_MUXInst_94_U1 ( .A(Red_Feedback[94]), .B(Red_Input[94]), 
        .S(rst), .Z(Red_MCInput[94]) );
  MUX2_X1 Red_InputMUX_MUXInst_95_U1 ( .A(Red_Feedback[95]), .B(Red_Input[95]), 
        .S(rst), .Z(Red_MCInput[95]) );
  MUX2_X1 Red_InputMUX_MUXInst_96_U1 ( .A(Red_Feedback[96]), .B(Red_Input[96]), 
        .S(rst), .Z(Red_MCInput[96]) );
  MUX2_X1 Red_InputMUX_MUXInst_97_U1 ( .A(Red_Feedback[97]), .B(Red_Input[97]), 
        .S(rst), .Z(Red_MCInput[97]) );
  MUX2_X1 Red_InputMUX_MUXInst_98_U1 ( .A(Red_Feedback[98]), .B(Red_Input[98]), 
        .S(rst), .Z(Red_MCInput[98]) );
  MUX2_X1 Red_InputMUX_MUXInst_99_U1 ( .A(Red_Feedback[99]), .B(Red_Input[99]), 
        .S(rst), .Z(Red_MCInput[99]) );
  MUX2_X1 Red_InputMUX_MUXInst_100_U1 ( .A(Red_Feedback[100]), .B(
        Red_Input[100]), .S(rst), .Z(Red_MCInput[100]) );
  MUX2_X1 Red_InputMUX_MUXInst_101_U1 ( .A(Red_Feedback[101]), .B(
        Red_Input[101]), .S(rst), .Z(Red_MCInput[101]) );
  MUX2_X1 Red_InputMUX_MUXInst_102_U1 ( .A(Red_Feedback[102]), .B(
        Red_Input[102]), .S(rst), .Z(Red_MCInput[102]) );
  MUX2_X1 Red_InputMUX_MUXInst_103_U1 ( .A(Red_Feedback[103]), .B(
        Red_Input[103]), .S(rst), .Z(Red_MCInput[103]) );
  MUX2_X1 Red_InputMUX_MUXInst_104_U1 ( .A(Red_Feedback[104]), .B(
        Red_Input[104]), .S(rst), .Z(Red_MCInput[104]) );
  MUX2_X1 Red_InputMUX_MUXInst_105_U1 ( .A(Red_Feedback[105]), .B(
        Red_Input[105]), .S(rst), .Z(Red_MCInput[105]) );
  MUX2_X1 Red_InputMUX_MUXInst_106_U1 ( .A(Red_Feedback[106]), .B(
        Red_Input[106]), .S(rst), .Z(Red_MCInput[106]) );
  MUX2_X1 Red_InputMUX_MUXInst_107_U1 ( .A(Red_Feedback[107]), .B(
        Red_Input[107]), .S(rst), .Z(Red_MCInput[107]) );
  MUX2_X1 Red_InputMUX_MUXInst_108_U1 ( .A(Red_Feedback[108]), .B(
        Red_Input[108]), .S(rst), .Z(Red_MCInput[108]) );
  MUX2_X1 Red_InputMUX_MUXInst_109_U1 ( .A(Red_Feedback[109]), .B(
        Red_Input[109]), .S(rst), .Z(Red_MCInput[109]) );
  MUX2_X1 Red_InputMUX_MUXInst_110_U1 ( .A(Red_Feedback[110]), .B(
        Red_Input[110]), .S(rst), .Z(Red_MCInput[110]) );
  MUX2_X1 Red_InputMUX_MUXInst_111_U1 ( .A(Red_Feedback[111]), .B(
        Red_Input[111]), .S(rst), .Z(Red_MCInput[111]) );
  XNOR2_X1 Red_MCInst_XOR_r0_Inst_0_U2 ( .A(Red_MCInst_XOR_r0_Inst_0_n5), .B(
        Red_MCOutput[28]), .ZN(Red_MCOutput[84]) );
  XNOR2_X1 Red_MCInst_XOR_r0_Inst_0_U1 ( .A(Red_MCOutput[0]), .B(
        Red_MCInput[84]), .ZN(Red_MCInst_XOR_r0_Inst_0_n5) );
  XOR2_X1 Red_MCInst_XOR_r1_Inst_0_U1 ( .A(Red_MCInput[56]), .B(
        Red_MCOutput[0]), .Z(Red_MCOutput[56]) );
  XNOR2_X1 Red_MCInst_XOR_r0_Inst_1_U2 ( .A(Red_MCInst_XOR_r0_Inst_1_n5), .B(
        Red_MCOutput[29]), .ZN(Red_MCOutput[85]) );
  XNOR2_X1 Red_MCInst_XOR_r0_Inst_1_U1 ( .A(Red_MCOutput[1]), .B(
        Red_MCInput[85]), .ZN(Red_MCInst_XOR_r0_Inst_1_n5) );
  XOR2_X1 Red_MCInst_XOR_r1_Inst_1_U1 ( .A(Red_MCInput[57]), .B(
        Red_MCOutput[1]), .Z(Red_MCOutput[57]) );
  XNOR2_X1 Red_MCInst_XOR_r0_Inst_2_U2 ( .A(Red_MCInst_XOR_r0_Inst_2_n5), .B(
        Red_MCOutput[30]), .ZN(Red_MCOutput[86]) );
  XNOR2_X1 Red_MCInst_XOR_r0_Inst_2_U1 ( .A(Red_MCOutput[2]), .B(
        Red_MCInput[86]), .ZN(Red_MCInst_XOR_r0_Inst_2_n5) );
  XOR2_X1 Red_MCInst_XOR_r1_Inst_2_U1 ( .A(Red_MCInput[58]), .B(
        Red_MCOutput[2]), .Z(Red_MCOutput[58]) );
  XNOR2_X1 Red_MCInst_XOR_r0_Inst_3_U2 ( .A(Red_MCInst_XOR_r0_Inst_3_n5), .B(
        Red_MCOutput[31]), .ZN(Red_MCOutput[87]) );
  XNOR2_X1 Red_MCInst_XOR_r0_Inst_3_U1 ( .A(Red_MCOutput[3]), .B(
        Red_MCInput[87]), .ZN(Red_MCInst_XOR_r0_Inst_3_n5) );
  XOR2_X1 Red_MCInst_XOR_r1_Inst_3_U1 ( .A(Red_MCInput[59]), .B(
        Red_MCOutput[3]), .Z(Red_MCOutput[59]) );
  XNOR2_X1 Red_MCInst_XOR_r0_Inst_4_U2 ( .A(Red_MCInst_XOR_r0_Inst_4_n5), .B(
        Red_MCOutput[32]), .ZN(Red_MCOutput[88]) );
  XNOR2_X1 Red_MCInst_XOR_r0_Inst_4_U1 ( .A(Red_MCOutput[4]), .B(
        Red_MCInput[88]), .ZN(Red_MCInst_XOR_r0_Inst_4_n5) );
  XOR2_X1 Red_MCInst_XOR_r1_Inst_4_U1 ( .A(Red_MCInput[60]), .B(
        Red_MCOutput[4]), .Z(Red_MCOutput[60]) );
  XNOR2_X1 Red_MCInst_XOR_r0_Inst_5_U2 ( .A(Red_MCInst_XOR_r0_Inst_5_n5), .B(
        Red_MCOutput[33]), .ZN(Red_MCOutput[89]) );
  XNOR2_X1 Red_MCInst_XOR_r0_Inst_5_U1 ( .A(Red_MCOutput[5]), .B(
        Red_MCInput[89]), .ZN(Red_MCInst_XOR_r0_Inst_5_n5) );
  XOR2_X1 Red_MCInst_XOR_r1_Inst_5_U1 ( .A(Red_MCInput[61]), .B(
        Red_MCOutput[5]), .Z(Red_MCOutput[61]) );
  XNOR2_X1 Red_MCInst_XOR_r0_Inst_6_U2 ( .A(Red_MCInst_XOR_r0_Inst_6_n5), .B(
        Red_MCOutput[34]), .ZN(Red_MCOutput[90]) );
  XNOR2_X1 Red_MCInst_XOR_r0_Inst_6_U1 ( .A(Red_MCOutput[6]), .B(
        Red_MCInput[90]), .ZN(Red_MCInst_XOR_r0_Inst_6_n5) );
  XOR2_X1 Red_MCInst_XOR_r1_Inst_6_U1 ( .A(Red_MCInput[62]), .B(
        Red_MCOutput[6]), .Z(Red_MCOutput[62]) );
  XNOR2_X1 Red_MCInst_XOR_r0_Inst_7_U2 ( .A(Red_MCInst_XOR_r0_Inst_7_n5), .B(
        Red_MCOutput[35]), .ZN(Red_MCOutput[91]) );
  XNOR2_X1 Red_MCInst_XOR_r0_Inst_7_U1 ( .A(Red_MCOutput[7]), .B(
        Red_MCInput[91]), .ZN(Red_MCInst_XOR_r0_Inst_7_n5) );
  XOR2_X1 Red_MCInst_XOR_r1_Inst_7_U1 ( .A(Red_MCInput[63]), .B(
        Red_MCOutput[7]), .Z(Red_MCOutput[63]) );
  XNOR2_X1 Red_MCInst_XOR_r0_Inst_8_U2 ( .A(Red_MCInst_XOR_r0_Inst_8_n5), .B(
        Red_MCOutput[36]), .ZN(Red_MCOutput[92]) );
  XNOR2_X1 Red_MCInst_XOR_r0_Inst_8_U1 ( .A(Red_MCOutput[8]), .B(
        Red_MCInput[92]), .ZN(Red_MCInst_XOR_r0_Inst_8_n5) );
  XOR2_X1 Red_MCInst_XOR_r1_Inst_8_U1 ( .A(Red_MCInput[64]), .B(
        Red_MCOutput[8]), .Z(Red_MCOutput[64]) );
  XNOR2_X1 Red_MCInst_XOR_r0_Inst_9_U2 ( .A(Red_MCInst_XOR_r0_Inst_9_n5), .B(
        Red_MCOutput[37]), .ZN(Red_MCOutput[93]) );
  XNOR2_X1 Red_MCInst_XOR_r0_Inst_9_U1 ( .A(Red_MCOutput[9]), .B(
        Red_MCInput[93]), .ZN(Red_MCInst_XOR_r0_Inst_9_n5) );
  XOR2_X1 Red_MCInst_XOR_r1_Inst_9_U1 ( .A(Red_MCInput[65]), .B(
        Red_MCOutput[9]), .Z(Red_MCOutput[65]) );
  XNOR2_X1 Red_MCInst_XOR_r0_Inst_10_U2 ( .A(Red_MCInst_XOR_r0_Inst_10_n5), 
        .B(Red_MCOutput[38]), .ZN(Red_MCOutput[94]) );
  XNOR2_X1 Red_MCInst_XOR_r0_Inst_10_U1 ( .A(Red_MCOutput[10]), .B(
        Red_MCInput[94]), .ZN(Red_MCInst_XOR_r0_Inst_10_n5) );
  XOR2_X1 Red_MCInst_XOR_r1_Inst_10_U1 ( .A(Red_MCInput[66]), .B(
        Red_MCOutput[10]), .Z(Red_MCOutput[66]) );
  XNOR2_X1 Red_MCInst_XOR_r0_Inst_11_U2 ( .A(Red_MCInst_XOR_r0_Inst_11_n5), 
        .B(Red_MCOutput[39]), .ZN(Red_MCOutput[95]) );
  XNOR2_X1 Red_MCInst_XOR_r0_Inst_11_U1 ( .A(Red_MCOutput[11]), .B(
        Red_MCInput[95]), .ZN(Red_MCInst_XOR_r0_Inst_11_n5) );
  XOR2_X1 Red_MCInst_XOR_r1_Inst_11_U1 ( .A(Red_MCInput[67]), .B(
        Red_MCOutput[11]), .Z(Red_MCOutput[67]) );
  XNOR2_X1 Red_MCInst_XOR_r0_Inst_12_U2 ( .A(Red_MCInst_XOR_r0_Inst_12_n5), 
        .B(Red_MCOutput[40]), .ZN(Red_MCOutput[96]) );
  XNOR2_X1 Red_MCInst_XOR_r0_Inst_12_U1 ( .A(Red_MCOutput[12]), .B(
        Red_MCInput[96]), .ZN(Red_MCInst_XOR_r0_Inst_12_n5) );
  XOR2_X1 Red_MCInst_XOR_r1_Inst_12_U1 ( .A(Red_MCInput[68]), .B(
        Red_MCOutput[12]), .Z(Red_MCOutput[68]) );
  XNOR2_X1 Red_MCInst_XOR_r0_Inst_13_U2 ( .A(Red_MCInst_XOR_r0_Inst_13_n5), 
        .B(Red_MCOutput[41]), .ZN(Red_MCOutput[97]) );
  XNOR2_X1 Red_MCInst_XOR_r0_Inst_13_U1 ( .A(Red_MCOutput[13]), .B(
        Red_MCInput[97]), .ZN(Red_MCInst_XOR_r0_Inst_13_n5) );
  XOR2_X1 Red_MCInst_XOR_r1_Inst_13_U1 ( .A(Red_MCInput[69]), .B(
        Red_MCOutput[13]), .Z(Red_MCOutput[69]) );
  XNOR2_X1 Red_MCInst_XOR_r0_Inst_14_U2 ( .A(Red_MCInst_XOR_r0_Inst_14_n5), 
        .B(Red_MCOutput[42]), .ZN(Red_MCOutput[98]) );
  XNOR2_X1 Red_MCInst_XOR_r0_Inst_14_U1 ( .A(Red_MCOutput[14]), .B(
        Red_MCInput[98]), .ZN(Red_MCInst_XOR_r0_Inst_14_n5) );
  XOR2_X1 Red_MCInst_XOR_r1_Inst_14_U1 ( .A(Red_MCInput[70]), .B(
        Red_MCOutput[14]), .Z(Red_MCOutput[70]) );
  XNOR2_X1 Red_MCInst_XOR_r0_Inst_15_U2 ( .A(Red_MCInst_XOR_r0_Inst_15_n5), 
        .B(Red_MCOutput[43]), .ZN(Red_MCOutput[99]) );
  XNOR2_X1 Red_MCInst_XOR_r0_Inst_15_U1 ( .A(Red_MCOutput[15]), .B(
        Red_MCInput[99]), .ZN(Red_MCInst_XOR_r0_Inst_15_n5) );
  XOR2_X1 Red_MCInst_XOR_r1_Inst_15_U1 ( .A(Red_MCInput[71]), .B(
        Red_MCOutput[15]), .Z(Red_MCOutput[71]) );
  XNOR2_X1 Red_MCInst_XOR_r0_Inst_16_U2 ( .A(Red_MCInst_XOR_r0_Inst_16_n5), 
        .B(Red_MCOutput[44]), .ZN(Red_MCOutput[100]) );
  XNOR2_X1 Red_MCInst_XOR_r0_Inst_16_U1 ( .A(Red_MCOutput[16]), .B(
        Red_MCInput[100]), .ZN(Red_MCInst_XOR_r0_Inst_16_n5) );
  XOR2_X1 Red_MCInst_XOR_r1_Inst_16_U1 ( .A(Red_MCInput[72]), .B(
        Red_MCOutput[16]), .Z(Red_MCOutput[72]) );
  XNOR2_X1 Red_MCInst_XOR_r0_Inst_17_U2 ( .A(Red_MCInst_XOR_r0_Inst_17_n5), 
        .B(Red_MCOutput[45]), .ZN(Red_MCOutput[101]) );
  XNOR2_X1 Red_MCInst_XOR_r0_Inst_17_U1 ( .A(Red_MCOutput[17]), .B(
        Red_MCInput[101]), .ZN(Red_MCInst_XOR_r0_Inst_17_n5) );
  XOR2_X1 Red_MCInst_XOR_r1_Inst_17_U1 ( .A(Red_MCInput[73]), .B(
        Red_MCOutput[17]), .Z(Red_MCOutput[73]) );
  XNOR2_X1 Red_MCInst_XOR_r0_Inst_18_U2 ( .A(Red_MCInst_XOR_r0_Inst_18_n5), 
        .B(Red_MCOutput[46]), .ZN(Red_MCOutput[102]) );
  XNOR2_X1 Red_MCInst_XOR_r0_Inst_18_U1 ( .A(Red_MCOutput[18]), .B(
        Red_MCInput[102]), .ZN(Red_MCInst_XOR_r0_Inst_18_n5) );
  XOR2_X1 Red_MCInst_XOR_r1_Inst_18_U1 ( .A(Red_MCInput[74]), .B(
        Red_MCOutput[18]), .Z(Red_MCOutput[74]) );
  XNOR2_X1 Red_MCInst_XOR_r0_Inst_19_U2 ( .A(Red_MCInst_XOR_r0_Inst_19_n5), 
        .B(Red_MCOutput[47]), .ZN(Red_MCOutput[103]) );
  XNOR2_X1 Red_MCInst_XOR_r0_Inst_19_U1 ( .A(Red_MCOutput[19]), .B(
        Red_MCInput[103]), .ZN(Red_MCInst_XOR_r0_Inst_19_n5) );
  XOR2_X1 Red_MCInst_XOR_r1_Inst_19_U1 ( .A(Red_MCInput[75]), .B(
        Red_MCOutput[19]), .Z(Red_MCOutput[75]) );
  XNOR2_X1 Red_MCInst_XOR_r0_Inst_20_U2 ( .A(Red_MCInst_XOR_r0_Inst_20_n5), 
        .B(Red_MCOutput[48]), .ZN(Red_MCOutput[104]) );
  XNOR2_X1 Red_MCInst_XOR_r0_Inst_20_U1 ( .A(Red_MCOutput[20]), .B(
        Red_MCInput[104]), .ZN(Red_MCInst_XOR_r0_Inst_20_n5) );
  XOR2_X1 Red_MCInst_XOR_r1_Inst_20_U1 ( .A(Red_MCInput[76]), .B(
        Red_MCOutput[20]), .Z(Red_MCOutput[76]) );
  XNOR2_X1 Red_MCInst_XOR_r0_Inst_21_U2 ( .A(Red_MCInst_XOR_r0_Inst_21_n5), 
        .B(Red_MCOutput[49]), .ZN(Red_MCOutput[105]) );
  XNOR2_X1 Red_MCInst_XOR_r0_Inst_21_U1 ( .A(Red_MCOutput[21]), .B(
        Red_MCInput[105]), .ZN(Red_MCInst_XOR_r0_Inst_21_n5) );
  XOR2_X1 Red_MCInst_XOR_r1_Inst_21_U1 ( .A(Red_MCInput[77]), .B(
        Red_MCOutput[21]), .Z(Red_MCOutput[77]) );
  XNOR2_X1 Red_MCInst_XOR_r0_Inst_22_U2 ( .A(Red_MCInst_XOR_r0_Inst_22_n5), 
        .B(Red_MCOutput[50]), .ZN(Red_MCOutput[106]) );
  XNOR2_X1 Red_MCInst_XOR_r0_Inst_22_U1 ( .A(Red_MCOutput[22]), .B(
        Red_MCInput[106]), .ZN(Red_MCInst_XOR_r0_Inst_22_n5) );
  XOR2_X1 Red_MCInst_XOR_r1_Inst_22_U1 ( .A(Red_MCInput[78]), .B(
        Red_MCOutput[22]), .Z(Red_MCOutput[78]) );
  XNOR2_X1 Red_MCInst_XOR_r0_Inst_23_U2 ( .A(Red_MCInst_XOR_r0_Inst_23_n5), 
        .B(Red_MCOutput[51]), .ZN(Red_MCOutput[107]) );
  XNOR2_X1 Red_MCInst_XOR_r0_Inst_23_U1 ( .A(Red_MCOutput[23]), .B(
        Red_MCInput[107]), .ZN(Red_MCInst_XOR_r0_Inst_23_n5) );
  XOR2_X1 Red_MCInst_XOR_r1_Inst_23_U1 ( .A(Red_MCInput[79]), .B(
        Red_MCOutput[23]), .Z(Red_MCOutput[79]) );
  XNOR2_X1 Red_MCInst_XOR_r0_Inst_24_U2 ( .A(Red_MCInst_XOR_r0_Inst_24_n5), 
        .B(Red_MCOutput[52]), .ZN(Red_MCOutput[108]) );
  XNOR2_X1 Red_MCInst_XOR_r0_Inst_24_U1 ( .A(Red_MCOutput[24]), .B(
        Red_MCInput[108]), .ZN(Red_MCInst_XOR_r0_Inst_24_n5) );
  XOR2_X1 Red_MCInst_XOR_r1_Inst_24_U1 ( .A(Red_MCInput[80]), .B(
        Red_MCOutput[24]), .Z(Red_MCOutput[80]) );
  XNOR2_X1 Red_MCInst_XOR_r0_Inst_25_U2 ( .A(Red_MCInst_XOR_r0_Inst_25_n5), 
        .B(Red_MCOutput[53]), .ZN(Red_MCOutput[109]) );
  XNOR2_X1 Red_MCInst_XOR_r0_Inst_25_U1 ( .A(Red_MCOutput[25]), .B(
        Red_MCInput[109]), .ZN(Red_MCInst_XOR_r0_Inst_25_n5) );
  XOR2_X1 Red_MCInst_XOR_r1_Inst_25_U1 ( .A(Red_MCInput[81]), .B(
        Red_MCOutput[25]), .Z(Red_MCOutput[81]) );
  XNOR2_X1 Red_MCInst_XOR_r0_Inst_26_U2 ( .A(Red_MCInst_XOR_r0_Inst_26_n5), 
        .B(Red_MCOutput[54]), .ZN(Red_MCOutput[110]) );
  XNOR2_X1 Red_MCInst_XOR_r0_Inst_26_U1 ( .A(Red_MCOutput[26]), .B(
        Red_MCInput[110]), .ZN(Red_MCInst_XOR_r0_Inst_26_n5) );
  XOR2_X1 Red_MCInst_XOR_r1_Inst_26_U1 ( .A(Red_MCInput[82]), .B(
        Red_MCOutput[26]), .Z(Red_MCOutput[82]) );
  XNOR2_X1 Red_MCInst_XOR_r0_Inst_27_U2 ( .A(Red_MCInst_XOR_r0_Inst_27_n5), 
        .B(Red_MCOutput[55]), .ZN(Red_MCOutput[111]) );
  XNOR2_X1 Red_MCInst_XOR_r0_Inst_27_U1 ( .A(Red_MCOutput[27]), .B(
        Red_MCInput[111]), .ZN(Red_MCInst_XOR_r0_Inst_27_n5) );
  XOR2_X1 Red_MCInst_XOR_r1_Inst_27_U1 ( .A(Red_MCInput[83]), .B(
        Red_MCOutput[27]), .Z(Red_MCOutput[83]) );
  XOR2_X1 Red_AddKeyXOR1_XORInst_0_0_U1 ( .A(Red_MCOutput[84]), .B(
        Red_SelectedKey[84]), .Z(Red_AddRoundKeyOutput[84]) );
  XOR2_X1 Red_AddKeyXOR1_XORInst_0_1_U1 ( .A(Red_MCOutput[85]), .B(
        Red_SelectedKey[85]), .Z(Red_AddRoundKeyOutput[85]) );
  XOR2_X1 Red_AddKeyXOR1_XORInst_0_2_U1 ( .A(Red_MCOutput[86]), .B(
        Red_SelectedKey[86]), .Z(Red_AddRoundKeyOutput[86]) );
  XOR2_X1 Red_AddKeyXOR1_XORInst_0_3_U1 ( .A(Red_MCOutput[87]), .B(
        Red_SelectedKey[87]), .Z(Red_AddRoundKeyOutput[87]) );
  XOR2_X1 Red_AddKeyXOR1_XORInst_0_4_U1 ( .A(Red_MCOutput[88]), .B(
        Red_SelectedKey[88]), .Z(Red_AddRoundKeyOutput[88]) );
  XOR2_X1 Red_AddKeyXOR1_XORInst_0_5_U1 ( .A(Red_MCOutput[89]), .B(
        Red_SelectedKey[89]), .Z(Red_AddRoundKeyOutput[89]) );
  XOR2_X1 Red_AddKeyXOR1_XORInst_0_6_U1 ( .A(Red_MCOutput[90]), .B(
        Red_SelectedKey[90]), .Z(Red_AddRoundKeyOutput[90]) );
  XOR2_X1 Red_AddKeyXOR1_XORInst_1_0_U1 ( .A(Red_MCOutput[91]), .B(
        Red_SelectedKey[91]), .Z(Red_AddRoundKeyOutput[91]) );
  XOR2_X1 Red_AddKeyXOR1_XORInst_1_1_U1 ( .A(Red_MCOutput[92]), .B(
        Red_SelectedKey[92]), .Z(Red_AddRoundKeyOutput[92]) );
  XOR2_X1 Red_AddKeyXOR1_XORInst_1_2_U1 ( .A(Red_MCOutput[93]), .B(
        Red_SelectedKey[93]), .Z(Red_AddRoundKeyOutput[93]) );
  XOR2_X1 Red_AddKeyXOR1_XORInst_1_3_U1 ( .A(Red_MCOutput[94]), .B(
        Red_SelectedKey[94]), .Z(Red_AddRoundKeyOutput[94]) );
  XOR2_X1 Red_AddKeyXOR1_XORInst_1_4_U1 ( .A(Red_MCOutput[95]), .B(
        Red_SelectedKey[95]), .Z(Red_AddRoundKeyOutput[95]) );
  XOR2_X1 Red_AddKeyXOR1_XORInst_1_5_U1 ( .A(Red_MCOutput[96]), .B(
        Red_SelectedKey[96]), .Z(Red_AddRoundKeyOutput[96]) );
  XOR2_X1 Red_AddKeyXOR1_XORInst_1_6_U1 ( .A(Red_MCOutput[97]), .B(
        Red_SelectedKey[97]), .Z(Red_AddRoundKeyOutput[97]) );
  XOR2_X1 Red_AddKeyXOR1_XORInst_2_0_U1 ( .A(Red_MCOutput[98]), .B(
        Red_SelectedKey[98]), .Z(Red_AddRoundKeyOutput[98]) );
  XOR2_X1 Red_AddKeyXOR1_XORInst_2_1_U1 ( .A(Red_MCOutput[99]), .B(
        Red_SelectedKey[99]), .Z(Red_AddRoundKeyOutput[99]) );
  XOR2_X1 Red_AddKeyXOR1_XORInst_2_2_U1 ( .A(Red_MCOutput[100]), .B(
        Red_SelectedKey[100]), .Z(Red_AddRoundKeyOutput[100]) );
  XOR2_X1 Red_AddKeyXOR1_XORInst_2_3_U1 ( .A(Red_MCOutput[101]), .B(
        Red_SelectedKey[101]), .Z(Red_AddRoundKeyOutput[101]) );
  XOR2_X1 Red_AddKeyXOR1_XORInst_2_4_U1 ( .A(Red_MCOutput[102]), .B(
        Red_SelectedKey[102]), .Z(Red_AddRoundKeyOutput[102]) );
  XOR2_X1 Red_AddKeyXOR1_XORInst_2_5_U1 ( .A(Red_MCOutput[103]), .B(
        Red_SelectedKey[103]), .Z(Red_AddRoundKeyOutput[103]) );
  XOR2_X1 Red_AddKeyXOR1_XORInst_2_6_U1 ( .A(Red_MCOutput[104]), .B(
        Red_SelectedKey[104]), .Z(Red_AddRoundKeyOutput[104]) );
  XOR2_X1 Red_AddKeyXOR1_XORInst_3_0_U1 ( .A(Red_MCOutput[105]), .B(
        Red_SelectedKey[105]), .Z(Red_AddRoundKeyOutput[105]) );
  XOR2_X1 Red_AddKeyXOR1_XORInst_3_1_U1 ( .A(Red_MCOutput[106]), .B(
        Red_SelectedKey[106]), .Z(Red_AddRoundKeyOutput[106]) );
  XOR2_X1 Red_AddKeyXOR1_XORInst_3_2_U1 ( .A(Red_MCOutput[107]), .B(
        Red_SelectedKey[107]), .Z(Red_AddRoundKeyOutput[107]) );
  XOR2_X1 Red_AddKeyXOR1_XORInst_3_3_U1 ( .A(Red_MCOutput[108]), .B(
        Red_SelectedKey[108]), .Z(Red_AddRoundKeyOutput[108]) );
  XOR2_X1 Red_AddKeyXOR1_XORInst_3_4_U1 ( .A(Red_MCOutput[109]), .B(
        Red_SelectedKey[109]), .Z(Red_AddRoundKeyOutput[109]) );
  XOR2_X1 Red_AddKeyXOR1_XORInst_3_5_U1 ( .A(Red_MCOutput[110]), .B(
        Red_SelectedKey[110]), .Z(Red_AddRoundKeyOutput[110]) );
  XOR2_X1 Red_AddKeyXOR1_XORInst_3_6_U1 ( .A(Red_MCOutput[111]), .B(
        Red_SelectedKey[111]), .Z(Red_AddRoundKeyOutput[111]) );
  XNOR2_X1 Red_AddKeyConstXOR_XORInst_0_0_U2 ( .A(
        Red_AddKeyConstXOR_XORInst_0_0_n5), .B(Red_SelectedKey[70]), .ZN(
        Red_AddRoundKeyOutput[70]) );
  XNOR2_X1 Red_AddKeyConstXOR_XORInst_0_0_U1 ( .A(Red_RoundConstant[0]), .B(
        Red_MCOutput[70]), .ZN(Red_AddKeyConstXOR_XORInst_0_0_n5) );
  XNOR2_X1 Red_AddKeyConstXOR_XORInst_0_1_U2 ( .A(
        Red_AddKeyConstXOR_XORInst_0_1_n5), .B(Red_SelectedKey[71]), .ZN(
        Red_AddRoundKeyOutput[71]) );
  XNOR2_X1 Red_AddKeyConstXOR_XORInst_0_1_U1 ( .A(Red_RoundConstant[1]), .B(
        Red_MCOutput[71]), .ZN(Red_AddKeyConstXOR_XORInst_0_1_n5) );
  XNOR2_X1 Red_AddKeyConstXOR_XORInst_0_2_U2 ( .A(
        Red_AddKeyConstXOR_XORInst_0_2_n5), .B(Red_SelectedKey[72]), .ZN(
        Red_AddRoundKeyOutput[72]) );
  XNOR2_X1 Red_AddKeyConstXOR_XORInst_0_2_U1 ( .A(Red_RoundConstant[2]), .B(
        Red_MCOutput[72]), .ZN(Red_AddKeyConstXOR_XORInst_0_2_n5) );
  XNOR2_X1 Red_AddKeyConstXOR_XORInst_0_3_U2 ( .A(
        Red_AddKeyConstXOR_XORInst_0_3_n5), .B(Red_SelectedKey[73]), .ZN(
        Red_AddRoundKeyOutput[73]) );
  XNOR2_X1 Red_AddKeyConstXOR_XORInst_0_3_U1 ( .A(Red_RoundConstant[3]), .B(
        Red_MCOutput[73]), .ZN(Red_AddKeyConstXOR_XORInst_0_3_n5) );
  XNOR2_X1 Red_AddKeyConstXOR_XORInst_0_4_U2 ( .A(
        Red_AddKeyConstXOR_XORInst_0_4_n5), .B(Red_SelectedKey[74]), .ZN(
        Red_AddRoundKeyOutput[74]) );
  XNOR2_X1 Red_AddKeyConstXOR_XORInst_0_4_U1 ( .A(Red_RoundConstant[4]), .B(
        Red_MCOutput[74]), .ZN(Red_AddKeyConstXOR_XORInst_0_4_n5) );
  XNOR2_X1 Red_AddKeyConstXOR_XORInst_0_5_U2 ( .A(
        Red_AddKeyConstXOR_XORInst_0_5_n5), .B(Red_SelectedKey[75]), .ZN(
        Red_AddRoundKeyOutput[75]) );
  XNOR2_X1 Red_AddKeyConstXOR_XORInst_0_5_U1 ( .A(Red_RoundConstant[5]), .B(
        Red_MCOutput[75]), .ZN(Red_AddKeyConstXOR_XORInst_0_5_n5) );
  XNOR2_X1 Red_AddKeyConstXOR_XORInst_0_6_U2 ( .A(
        Red_AddKeyConstXOR_XORInst_0_6_n5), .B(Red_SelectedKey[76]), .ZN(
        Red_AddRoundKeyOutput[76]) );
  XNOR2_X1 Red_AddKeyConstXOR_XORInst_0_6_U1 ( .A(Red_RoundConstant[6]), .B(
        Red_MCOutput[76]), .ZN(Red_AddKeyConstXOR_XORInst_0_6_n5) );
  XNOR2_X1 Red_AddKeyConstXOR_XORInst_1_0_U2 ( .A(
        Red_AddKeyConstXOR_XORInst_1_0_n5), .B(Red_SelectedKey[77]), .ZN(
        Red_AddRoundKeyOutput[77]) );
  XNOR2_X1 Red_AddKeyConstXOR_XORInst_1_0_U1 ( .A(Red_RoundConstant[7]), .B(
        Red_MCOutput[77]), .ZN(Red_AddKeyConstXOR_XORInst_1_0_n5) );
  XNOR2_X1 Red_AddKeyConstXOR_XORInst_1_1_U2 ( .A(
        Red_AddKeyConstXOR_XORInst_1_1_n5), .B(Red_SelectedKey[78]), .ZN(
        Red_AddRoundKeyOutput[78]) );
  XNOR2_X1 Red_AddKeyConstXOR_XORInst_1_1_U1 ( .A(Red_RoundConstant[8]), .B(
        Red_MCOutput[78]), .ZN(Red_AddKeyConstXOR_XORInst_1_1_n5) );
  XNOR2_X1 Red_AddKeyConstXOR_XORInst_1_2_U2 ( .A(
        Red_AddKeyConstXOR_XORInst_1_2_n5), .B(Red_SelectedKey[79]), .ZN(
        Red_AddRoundKeyOutput[79]) );
  XNOR2_X1 Red_AddKeyConstXOR_XORInst_1_2_U1 ( .A(Red_RoundConstant[9]), .B(
        Red_MCOutput[79]), .ZN(Red_AddKeyConstXOR_XORInst_1_2_n5) );
  XNOR2_X1 Red_AddKeyConstXOR_XORInst_1_3_U2 ( .A(
        Red_AddKeyConstXOR_XORInst_1_3_n5), .B(Red_SelectedKey[80]), .ZN(
        Red_AddRoundKeyOutput[80]) );
  XNOR2_X1 Red_AddKeyConstXOR_XORInst_1_3_U1 ( .A(Red_RoundConstant[10]), .B(
        Red_MCOutput[80]), .ZN(Red_AddKeyConstXOR_XORInst_1_3_n5) );
  XNOR2_X1 Red_AddKeyConstXOR_XORInst_1_4_U2 ( .A(
        Red_AddKeyConstXOR_XORInst_1_4_n5), .B(Red_SelectedKey[81]), .ZN(
        Red_AddRoundKeyOutput[81]) );
  XNOR2_X1 Red_AddKeyConstXOR_XORInst_1_4_U1 ( .A(Red_RoundConstant[11]), .B(
        Red_MCOutput[81]), .ZN(Red_AddKeyConstXOR_XORInst_1_4_n5) );
  XNOR2_X1 Red_AddKeyConstXOR_XORInst_1_5_U2 ( .A(
        Red_AddKeyConstXOR_XORInst_1_5_n5), .B(Red_SelectedKey[82]), .ZN(
        Red_AddRoundKeyOutput[82]) );
  XNOR2_X1 Red_AddKeyConstXOR_XORInst_1_5_U1 ( .A(Red_RoundConstant[12]), .B(
        Red_MCOutput[82]), .ZN(Red_AddKeyConstXOR_XORInst_1_5_n5) );
  XNOR2_X1 Red_AddKeyConstXOR_XORInst_1_6_U2 ( .A(
        Red_AddKeyConstXOR_XORInst_1_6_n5), .B(Red_SelectedKey[83]), .ZN(
        Red_AddRoundKeyOutput[83]) );
  XNOR2_X1 Red_AddKeyConstXOR_XORInst_1_6_U1 ( .A(Red_RoundConstant[13]), .B(
        Red_MCOutput[83]), .ZN(Red_AddKeyConstXOR_XORInst_1_6_n5) );
  XOR2_X1 Red_AddKeyXOR2_XORInst_0_0_U1 ( .A(Red_MCOutput[0]), .B(
        Red_SelectedKey[0]), .Z(Red_AddRoundKeyOutput[0]) );
  XOR2_X1 Red_AddKeyXOR2_XORInst_0_1_U1 ( .A(Red_MCOutput[1]), .B(
        Red_SelectedKey[1]), .Z(Red_AddRoundKeyOutput[1]) );
  XOR2_X1 Red_AddKeyXOR2_XORInst_0_2_U1 ( .A(Red_MCOutput[2]), .B(
        Red_SelectedKey[2]), .Z(Red_AddRoundKeyOutput[2]) );
  XOR2_X1 Red_AddKeyXOR2_XORInst_0_3_U1 ( .A(Red_MCOutput[3]), .B(
        Red_SelectedKey[3]), .Z(Red_AddRoundKeyOutput[3]) );
  XOR2_X1 Red_AddKeyXOR2_XORInst_0_4_U1 ( .A(Red_MCOutput[4]), .B(
        Red_SelectedKey[4]), .Z(Red_AddRoundKeyOutput[4]) );
  XOR2_X1 Red_AddKeyXOR2_XORInst_0_5_U1 ( .A(Red_MCOutput[5]), .B(
        Red_SelectedKey[5]), .Z(Red_AddRoundKeyOutput[5]) );
  XOR2_X1 Red_AddKeyXOR2_XORInst_0_6_U1 ( .A(Red_MCOutput[6]), .B(
        Red_SelectedKey[6]), .Z(Red_AddRoundKeyOutput[6]) );
  XOR2_X1 Red_AddKeyXOR2_XORInst_1_0_U1 ( .A(Red_MCOutput[7]), .B(
        Red_SelectedKey[7]), .Z(Red_AddRoundKeyOutput[7]) );
  XOR2_X1 Red_AddKeyXOR2_XORInst_1_1_U1 ( .A(Red_MCOutput[8]), .B(
        Red_SelectedKey[8]), .Z(Red_AddRoundKeyOutput[8]) );
  XOR2_X1 Red_AddKeyXOR2_XORInst_1_2_U1 ( .A(Red_MCOutput[9]), .B(
        Red_SelectedKey[9]), .Z(Red_AddRoundKeyOutput[9]) );
  XOR2_X1 Red_AddKeyXOR2_XORInst_1_3_U1 ( .A(Red_MCOutput[10]), .B(
        Red_SelectedKey[10]), .Z(Red_AddRoundKeyOutput[10]) );
  XOR2_X1 Red_AddKeyXOR2_XORInst_1_4_U1 ( .A(Red_MCOutput[11]), .B(
        Red_SelectedKey[11]), .Z(Red_AddRoundKeyOutput[11]) );
  XOR2_X1 Red_AddKeyXOR2_XORInst_1_5_U1 ( .A(Red_MCOutput[12]), .B(
        Red_SelectedKey[12]), .Z(Red_AddRoundKeyOutput[12]) );
  XOR2_X1 Red_AddKeyXOR2_XORInst_1_6_U1 ( .A(Red_MCOutput[13]), .B(
        Red_SelectedKey[13]), .Z(Red_AddRoundKeyOutput[13]) );
  XOR2_X1 Red_AddKeyXOR2_XORInst_2_0_U1 ( .A(Red_MCOutput[14]), .B(
        Red_SelectedKey[14]), .Z(Red_AddRoundKeyOutput[14]) );
  XOR2_X1 Red_AddKeyXOR2_XORInst_2_1_U1 ( .A(Red_MCOutput[15]), .B(
        Red_SelectedKey[15]), .Z(Red_AddRoundKeyOutput[15]) );
  XOR2_X1 Red_AddKeyXOR2_XORInst_2_2_U1 ( .A(Red_MCOutput[16]), .B(
        Red_SelectedKey[16]), .Z(Red_AddRoundKeyOutput[16]) );
  XOR2_X1 Red_AddKeyXOR2_XORInst_2_3_U1 ( .A(Red_MCOutput[17]), .B(
        Red_SelectedKey[17]), .Z(Red_AddRoundKeyOutput[17]) );
  XOR2_X1 Red_AddKeyXOR2_XORInst_2_4_U1 ( .A(Red_MCOutput[18]), .B(
        Red_SelectedKey[18]), .Z(Red_AddRoundKeyOutput[18]) );
  XOR2_X1 Red_AddKeyXOR2_XORInst_2_5_U1 ( .A(Red_MCOutput[19]), .B(
        Red_SelectedKey[19]), .Z(Red_AddRoundKeyOutput[19]) );
  XOR2_X1 Red_AddKeyXOR2_XORInst_2_6_U1 ( .A(Red_MCOutput[20]), .B(
        Red_SelectedKey[20]), .Z(Red_AddRoundKeyOutput[20]) );
  XOR2_X1 Red_AddKeyXOR2_XORInst_3_0_U1 ( .A(Red_MCOutput[21]), .B(
        Red_SelectedKey[21]), .Z(Red_AddRoundKeyOutput[21]) );
  XOR2_X1 Red_AddKeyXOR2_XORInst_3_1_U1 ( .A(Red_MCOutput[22]), .B(
        Red_SelectedKey[22]), .Z(Red_AddRoundKeyOutput[22]) );
  XOR2_X1 Red_AddKeyXOR2_XORInst_3_2_U1 ( .A(Red_MCOutput[23]), .B(
        Red_SelectedKey[23]), .Z(Red_AddRoundKeyOutput[23]) );
  XOR2_X1 Red_AddKeyXOR2_XORInst_3_3_U1 ( .A(Red_MCOutput[24]), .B(
        Red_SelectedKey[24]), .Z(Red_AddRoundKeyOutput[24]) );
  XOR2_X1 Red_AddKeyXOR2_XORInst_3_4_U1 ( .A(Red_MCOutput[25]), .B(
        Red_SelectedKey[25]), .Z(Red_AddRoundKeyOutput[25]) );
  XOR2_X1 Red_AddKeyXOR2_XORInst_3_5_U1 ( .A(Red_MCOutput[26]), .B(
        Red_SelectedKey[26]), .Z(Red_AddRoundKeyOutput[26]) );
  XOR2_X1 Red_AddKeyXOR2_XORInst_3_6_U1 ( .A(Red_MCOutput[27]), .B(
        Red_SelectedKey[27]), .Z(Red_AddRoundKeyOutput[27]) );
  XOR2_X1 Red_AddKeyXOR2_XORInst_4_0_U1 ( .A(Red_MCOutput[28]), .B(
        Red_SelectedKey[28]), .Z(Red_AddRoundKeyOutput[28]) );
  XOR2_X1 Red_AddKeyXOR2_XORInst_4_1_U1 ( .A(Red_MCOutput[29]), .B(
        Red_SelectedKey[29]), .Z(Red_AddRoundKeyOutput[29]) );
  XOR2_X1 Red_AddKeyXOR2_XORInst_4_2_U1 ( .A(Red_MCOutput[30]), .B(
        Red_SelectedKey[30]), .Z(Red_AddRoundKeyOutput[30]) );
  XOR2_X1 Red_AddKeyXOR2_XORInst_4_3_U1 ( .A(Red_MCOutput[31]), .B(
        Red_SelectedKey[31]), .Z(Red_AddRoundKeyOutput[31]) );
  XOR2_X1 Red_AddKeyXOR2_XORInst_4_4_U1 ( .A(Red_MCOutput[32]), .B(
        Red_SelectedKey[32]), .Z(Red_AddRoundKeyOutput[32]) );
  XOR2_X1 Red_AddKeyXOR2_XORInst_4_5_U1 ( .A(Red_MCOutput[33]), .B(
        Red_SelectedKey[33]), .Z(Red_AddRoundKeyOutput[33]) );
  XOR2_X1 Red_AddKeyXOR2_XORInst_4_6_U1 ( .A(Red_MCOutput[34]), .B(
        Red_SelectedKey[34]), .Z(Red_AddRoundKeyOutput[34]) );
  XOR2_X1 Red_AddKeyXOR2_XORInst_5_0_U1 ( .A(Red_MCOutput[35]), .B(
        Red_SelectedKey[35]), .Z(Red_AddRoundKeyOutput[35]) );
  XOR2_X1 Red_AddKeyXOR2_XORInst_5_1_U1 ( .A(Red_MCOutput[36]), .B(
        Red_SelectedKey[36]), .Z(Red_AddRoundKeyOutput[36]) );
  XOR2_X1 Red_AddKeyXOR2_XORInst_5_2_U1 ( .A(Red_MCOutput[37]), .B(
        Red_SelectedKey[37]), .Z(Red_AddRoundKeyOutput[37]) );
  XOR2_X1 Red_AddKeyXOR2_XORInst_5_3_U1 ( .A(Red_MCOutput[38]), .B(
        Red_SelectedKey[38]), .Z(Red_AddRoundKeyOutput[38]) );
  XOR2_X1 Red_AddKeyXOR2_XORInst_5_4_U1 ( .A(Red_MCOutput[39]), .B(
        Red_SelectedKey[39]), .Z(Red_AddRoundKeyOutput[39]) );
  XOR2_X1 Red_AddKeyXOR2_XORInst_5_5_U1 ( .A(Red_MCOutput[40]), .B(
        Red_SelectedKey[40]), .Z(Red_AddRoundKeyOutput[40]) );
  XOR2_X1 Red_AddKeyXOR2_XORInst_5_6_U1 ( .A(Red_MCOutput[41]), .B(
        Red_SelectedKey[41]), .Z(Red_AddRoundKeyOutput[41]) );
  XOR2_X1 Red_AddKeyXOR2_XORInst_6_0_U1 ( .A(Red_MCOutput[42]), .B(
        Red_SelectedKey[42]), .Z(Red_AddRoundKeyOutput[42]) );
  XOR2_X1 Red_AddKeyXOR2_XORInst_6_1_U1 ( .A(Red_MCOutput[43]), .B(
        Red_SelectedKey[43]), .Z(Red_AddRoundKeyOutput[43]) );
  XOR2_X1 Red_AddKeyXOR2_XORInst_6_2_U1 ( .A(Red_MCOutput[44]), .B(
        Red_SelectedKey[44]), .Z(Red_AddRoundKeyOutput[44]) );
  XOR2_X1 Red_AddKeyXOR2_XORInst_6_3_U1 ( .A(Red_MCOutput[45]), .B(
        Red_SelectedKey[45]), .Z(Red_AddRoundKeyOutput[45]) );
  XOR2_X1 Red_AddKeyXOR2_XORInst_6_4_U1 ( .A(Red_MCOutput[46]), .B(
        Red_SelectedKey[46]), .Z(Red_AddRoundKeyOutput[46]) );
  XOR2_X1 Red_AddKeyXOR2_XORInst_6_5_U1 ( .A(Red_MCOutput[47]), .B(
        Red_SelectedKey[47]), .Z(Red_AddRoundKeyOutput[47]) );
  XOR2_X1 Red_AddKeyXOR2_XORInst_6_6_U1 ( .A(Red_MCOutput[48]), .B(
        Red_SelectedKey[48]), .Z(Red_AddRoundKeyOutput[48]) );
  XOR2_X1 Red_AddKeyXOR2_XORInst_7_0_U1 ( .A(Red_MCOutput[49]), .B(
        Red_SelectedKey[49]), .Z(Red_AddRoundKeyOutput[49]) );
  XOR2_X1 Red_AddKeyXOR2_XORInst_7_1_U1 ( .A(Red_MCOutput[50]), .B(
        Red_SelectedKey[50]), .Z(Red_AddRoundKeyOutput[50]) );
  XOR2_X1 Red_AddKeyXOR2_XORInst_7_2_U1 ( .A(Red_MCOutput[51]), .B(
        Red_SelectedKey[51]), .Z(Red_AddRoundKeyOutput[51]) );
  XOR2_X1 Red_AddKeyXOR2_XORInst_7_3_U1 ( .A(Red_MCOutput[52]), .B(
        Red_SelectedKey[52]), .Z(Red_AddRoundKeyOutput[52]) );
  XOR2_X1 Red_AddKeyXOR2_XORInst_7_4_U1 ( .A(Red_MCOutput[53]), .B(
        Red_SelectedKey[53]), .Z(Red_AddRoundKeyOutput[53]) );
  XOR2_X1 Red_AddKeyXOR2_XORInst_7_5_U1 ( .A(Red_MCOutput[54]), .B(
        Red_SelectedKey[54]), .Z(Red_AddRoundKeyOutput[54]) );
  XOR2_X1 Red_AddKeyXOR2_XORInst_7_6_U1 ( .A(Red_MCOutput[55]), .B(
        Red_SelectedKey[55]), .Z(Red_AddRoundKeyOutput[55]) );
  XOR2_X1 Red_AddKeyXOR2_XORInst_8_0_U1 ( .A(Red_MCOutput[56]), .B(
        Red_SelectedKey[56]), .Z(Red_AddRoundKeyOutput[56]) );
  XOR2_X1 Red_AddKeyXOR2_XORInst_8_1_U1 ( .A(Red_MCOutput[57]), .B(
        Red_SelectedKey[57]), .Z(Red_AddRoundKeyOutput[57]) );
  XOR2_X1 Red_AddKeyXOR2_XORInst_8_2_U1 ( .A(Red_MCOutput[58]), .B(
        Red_SelectedKey[58]), .Z(Red_AddRoundKeyOutput[58]) );
  XOR2_X1 Red_AddKeyXOR2_XORInst_8_3_U1 ( .A(Red_MCOutput[59]), .B(
        Red_SelectedKey[59]), .Z(Red_AddRoundKeyOutput[59]) );
  XOR2_X1 Red_AddKeyXOR2_XORInst_8_4_U1 ( .A(Red_MCOutput[60]), .B(
        Red_SelectedKey[60]), .Z(Red_AddRoundKeyOutput[60]) );
  XOR2_X1 Red_AddKeyXOR2_XORInst_8_5_U1 ( .A(Red_MCOutput[61]), .B(
        Red_SelectedKey[61]), .Z(Red_AddRoundKeyOutput[61]) );
  XOR2_X1 Red_AddKeyXOR2_XORInst_8_6_U1 ( .A(Red_MCOutput[62]), .B(
        Red_SelectedKey[62]), .Z(Red_AddRoundKeyOutput[62]) );
  XOR2_X1 Red_AddKeyXOR2_XORInst_9_0_U1 ( .A(Red_MCOutput[63]), .B(
        Red_SelectedKey[63]), .Z(Red_AddRoundKeyOutput[63]) );
  XOR2_X1 Red_AddKeyXOR2_XORInst_9_1_U1 ( .A(Red_MCOutput[64]), .B(
        Red_SelectedKey[64]), .Z(Red_AddRoundKeyOutput[64]) );
  XOR2_X1 Red_AddKeyXOR2_XORInst_9_2_U1 ( .A(Red_MCOutput[65]), .B(
        Red_SelectedKey[65]), .Z(Red_AddRoundKeyOutput[65]) );
  XOR2_X1 Red_AddKeyXOR2_XORInst_9_3_U1 ( .A(Red_MCOutput[66]), .B(
        Red_SelectedKey[66]), .Z(Red_AddRoundKeyOutput[66]) );
  XOR2_X1 Red_AddKeyXOR2_XORInst_9_4_U1 ( .A(Red_MCOutput[67]), .B(
        Red_SelectedKey[67]), .Z(Red_AddRoundKeyOutput[67]) );
  XOR2_X1 Red_AddKeyXOR2_XORInst_9_5_U1 ( .A(Red_MCOutput[68]), .B(
        Red_SelectedKey[68]), .Z(Red_AddRoundKeyOutput[68]) );
  XOR2_X1 Red_AddKeyXOR2_XORInst_9_6_U1 ( .A(Red_MCOutput[69]), .B(
        Red_SelectedKey[69]), .Z(Red_AddRoundKeyOutput[69]) );
  DFF_X1 Red_StateReg_s_current_state_reg_0_ ( .D(Red_AddRoundKeyOutput[0]), 
        .CK(clk), .Q(Red_StateRegOutput[0]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_1_ ( .D(Red_AddRoundKeyOutput[1]), 
        .CK(clk), .Q(Red_StateRegOutput[1]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_2_ ( .D(Red_AddRoundKeyOutput[2]), 
        .CK(clk), .Q(Red_StateRegOutput[2]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_3_ ( .D(Red_AddRoundKeyOutput[3]), 
        .CK(clk), .Q(Red_StateRegOutput[3]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_4_ ( .D(Red_AddRoundKeyOutput[4]), 
        .CK(clk), .Q(Red_StateRegOutput[4]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_5_ ( .D(Red_AddRoundKeyOutput[5]), 
        .CK(clk), .Q(Red_StateRegOutput[5]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_6_ ( .D(Red_AddRoundKeyOutput[6]), 
        .CK(clk), .Q(Red_StateRegOutput[6]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_7_ ( .D(Red_AddRoundKeyOutput[7]), 
        .CK(clk), .Q(Red_StateRegOutput[7]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_8_ ( .D(Red_AddRoundKeyOutput[8]), 
        .CK(clk), .Q(Red_StateRegOutput[8]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_9_ ( .D(Red_AddRoundKeyOutput[9]), 
        .CK(clk), .Q(Red_StateRegOutput[9]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_10_ ( .D(Red_AddRoundKeyOutput[10]), 
        .CK(clk), .Q(Red_StateRegOutput[10]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_11_ ( .D(Red_AddRoundKeyOutput[11]), 
        .CK(clk), .Q(Red_StateRegOutput[11]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_12_ ( .D(Red_AddRoundKeyOutput[12]), 
        .CK(clk), .Q(Red_StateRegOutput[12]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_13_ ( .D(Red_AddRoundKeyOutput[13]), 
        .CK(clk), .Q(Red_StateRegOutput[13]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_14_ ( .D(Red_AddRoundKeyOutput[14]), 
        .CK(clk), .Q(Red_StateRegOutput[14]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_15_ ( .D(Red_AddRoundKeyOutput[15]), 
        .CK(clk), .Q(Red_StateRegOutput[15]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_16_ ( .D(Red_AddRoundKeyOutput[16]), 
        .CK(clk), .Q(Red_StateRegOutput[16]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_17_ ( .D(Red_AddRoundKeyOutput[17]), 
        .CK(clk), .Q(Red_StateRegOutput[17]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_18_ ( .D(Red_AddRoundKeyOutput[18]), 
        .CK(clk), .Q(Red_StateRegOutput[18]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_19_ ( .D(Red_AddRoundKeyOutput[19]), 
        .CK(clk), .Q(Red_StateRegOutput[19]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_20_ ( .D(Red_AddRoundKeyOutput[20]), 
        .CK(clk), .Q(Red_StateRegOutput[20]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_21_ ( .D(Red_AddRoundKeyOutput[21]), 
        .CK(clk), .Q(Red_StateRegOutput[21]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_22_ ( .D(Red_AddRoundKeyOutput[22]), 
        .CK(clk), .Q(Red_StateRegOutput[22]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_23_ ( .D(Red_AddRoundKeyOutput[23]), 
        .CK(clk), .Q(Red_StateRegOutput[23]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_24_ ( .D(Red_AddRoundKeyOutput[24]), 
        .CK(clk), .Q(Red_StateRegOutput[24]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_25_ ( .D(Red_AddRoundKeyOutput[25]), 
        .CK(clk), .Q(Red_StateRegOutput[25]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_26_ ( .D(Red_AddRoundKeyOutput[26]), 
        .CK(clk), .Q(Red_StateRegOutput[26]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_27_ ( .D(Red_AddRoundKeyOutput[27]), 
        .CK(clk), .Q(Red_StateRegOutput[27]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_28_ ( .D(Red_AddRoundKeyOutput[28]), 
        .CK(clk), .Q(Red_StateRegOutput[28]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_29_ ( .D(Red_AddRoundKeyOutput[29]), 
        .CK(clk), .Q(Red_StateRegOutput[29]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_30_ ( .D(Red_AddRoundKeyOutput[30]), 
        .CK(clk), .Q(Red_StateRegOutput[30]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_31_ ( .D(Red_AddRoundKeyOutput[31]), 
        .CK(clk), .Q(Red_StateRegOutput[31]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_32_ ( .D(Red_AddRoundKeyOutput[32]), 
        .CK(clk), .Q(Red_StateRegOutput[32]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_33_ ( .D(Red_AddRoundKeyOutput[33]), 
        .CK(clk), .Q(Red_StateRegOutput[33]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_34_ ( .D(Red_AddRoundKeyOutput[34]), 
        .CK(clk), .Q(Red_StateRegOutput[34]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_35_ ( .D(Red_AddRoundKeyOutput[35]), 
        .CK(clk), .Q(Red_StateRegOutput[35]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_36_ ( .D(Red_AddRoundKeyOutput[36]), 
        .CK(clk), .Q(Red_StateRegOutput[36]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_37_ ( .D(Red_AddRoundKeyOutput[37]), 
        .CK(clk), .Q(Red_StateRegOutput[37]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_38_ ( .D(Red_AddRoundKeyOutput[38]), 
        .CK(clk), .Q(Red_StateRegOutput[38]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_39_ ( .D(Red_AddRoundKeyOutput[39]), 
        .CK(clk), .Q(Red_StateRegOutput[39]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_40_ ( .D(Red_AddRoundKeyOutput[40]), 
        .CK(clk), .Q(Red_StateRegOutput[40]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_41_ ( .D(Red_AddRoundKeyOutput[41]), 
        .CK(clk), .Q(Red_StateRegOutput[41]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_42_ ( .D(Red_AddRoundKeyOutput[42]), 
        .CK(clk), .Q(Red_StateRegOutput[42]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_43_ ( .D(Red_AddRoundKeyOutput[43]), 
        .CK(clk), .Q(Red_StateRegOutput[43]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_44_ ( .D(Red_AddRoundKeyOutput[44]), 
        .CK(clk), .Q(Red_StateRegOutput[44]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_45_ ( .D(Red_AddRoundKeyOutput[45]), 
        .CK(clk), .Q(Red_StateRegOutput[45]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_46_ ( .D(Red_AddRoundKeyOutput[46]), 
        .CK(clk), .Q(Red_StateRegOutput[46]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_47_ ( .D(Red_AddRoundKeyOutput[47]), 
        .CK(clk), .Q(Red_StateRegOutput[47]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_48_ ( .D(Red_AddRoundKeyOutput[48]), 
        .CK(clk), .Q(Red_StateRegOutput[48]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_49_ ( .D(Red_AddRoundKeyOutput[49]), 
        .CK(clk), .Q(Red_StateRegOutput[49]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_50_ ( .D(Red_AddRoundKeyOutput[50]), 
        .CK(clk), .Q(Red_StateRegOutput[50]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_51_ ( .D(Red_AddRoundKeyOutput[51]), 
        .CK(clk), .Q(Red_StateRegOutput[51]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_52_ ( .D(Red_AddRoundKeyOutput[52]), 
        .CK(clk), .Q(Red_StateRegOutput[52]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_53_ ( .D(Red_AddRoundKeyOutput[53]), 
        .CK(clk), .Q(Red_StateRegOutput[53]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_54_ ( .D(Red_AddRoundKeyOutput[54]), 
        .CK(clk), .Q(Red_StateRegOutput[54]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_55_ ( .D(Red_AddRoundKeyOutput[55]), 
        .CK(clk), .Q(Red_StateRegOutput[55]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_56_ ( .D(Red_AddRoundKeyOutput[56]), 
        .CK(clk), .Q(Red_StateRegOutput[56]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_57_ ( .D(Red_AddRoundKeyOutput[57]), 
        .CK(clk), .Q(Red_StateRegOutput[57]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_58_ ( .D(Red_AddRoundKeyOutput[58]), 
        .CK(clk), .Q(Red_StateRegOutput[58]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_59_ ( .D(Red_AddRoundKeyOutput[59]), 
        .CK(clk), .Q(Red_StateRegOutput[59]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_60_ ( .D(Red_AddRoundKeyOutput[60]), 
        .CK(clk), .Q(Red_StateRegOutput[60]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_61_ ( .D(Red_AddRoundKeyOutput[61]), 
        .CK(clk), .Q(Red_StateRegOutput[61]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_62_ ( .D(Red_AddRoundKeyOutput[62]), 
        .CK(clk), .Q(Red_StateRegOutput[62]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_63_ ( .D(Red_AddRoundKeyOutput[63]), 
        .CK(clk), .Q(Red_StateRegOutput[63]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_64_ ( .D(Red_AddRoundKeyOutput[64]), 
        .CK(clk), .Q(Red_StateRegOutput[64]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_65_ ( .D(Red_AddRoundKeyOutput[65]), 
        .CK(clk), .Q(Red_StateRegOutput[65]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_66_ ( .D(Red_AddRoundKeyOutput[66]), 
        .CK(clk), .Q(Red_StateRegOutput[66]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_67_ ( .D(Red_AddRoundKeyOutput[67]), 
        .CK(clk), .Q(Red_StateRegOutput[67]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_68_ ( .D(Red_AddRoundKeyOutput[68]), 
        .CK(clk), .Q(Red_StateRegOutput[68]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_69_ ( .D(Red_AddRoundKeyOutput[69]), 
        .CK(clk), .Q(Red_StateRegOutput[69]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_70_ ( .D(Red_AddRoundKeyOutput[70]), 
        .CK(clk), .Q(Red_StateRegOutput[70]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_71_ ( .D(Red_AddRoundKeyOutput[71]), 
        .CK(clk), .Q(Red_StateRegOutput[71]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_72_ ( .D(Red_AddRoundKeyOutput[72]), 
        .CK(clk), .Q(Red_StateRegOutput[72]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_73_ ( .D(Red_AddRoundKeyOutput[73]), 
        .CK(clk), .Q(Red_StateRegOutput[73]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_74_ ( .D(Red_AddRoundKeyOutput[74]), 
        .CK(clk), .Q(Red_StateRegOutput[74]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_75_ ( .D(Red_AddRoundKeyOutput[75]), 
        .CK(clk), .Q(Red_StateRegOutput[75]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_76_ ( .D(Red_AddRoundKeyOutput[76]), 
        .CK(clk), .Q(Red_StateRegOutput[76]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_77_ ( .D(Red_AddRoundKeyOutput[77]), 
        .CK(clk), .Q(Red_StateRegOutput[77]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_78_ ( .D(Red_AddRoundKeyOutput[78]), 
        .CK(clk), .Q(Red_StateRegOutput[78]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_79_ ( .D(Red_AddRoundKeyOutput[79]), 
        .CK(clk), .Q(Red_StateRegOutput[79]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_80_ ( .D(Red_AddRoundKeyOutput[80]), 
        .CK(clk), .Q(Red_StateRegOutput[80]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_81_ ( .D(Red_AddRoundKeyOutput[81]), 
        .CK(clk), .Q(Red_StateRegOutput[81]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_82_ ( .D(Red_AddRoundKeyOutput[82]), 
        .CK(clk), .Q(Red_StateRegOutput[82]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_83_ ( .D(Red_AddRoundKeyOutput[83]), 
        .CK(clk), .Q(Red_StateRegOutput[83]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_84_ ( .D(Red_AddRoundKeyOutput[84]), 
        .CK(clk), .Q(Red_StateRegOutput[84]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_85_ ( .D(Red_AddRoundKeyOutput[85]), 
        .CK(clk), .Q(Red_StateRegOutput[85]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_86_ ( .D(Red_AddRoundKeyOutput[86]), 
        .CK(clk), .Q(Red_StateRegOutput[86]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_87_ ( .D(Red_AddRoundKeyOutput[87]), 
        .CK(clk), .Q(Red_StateRegOutput[87]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_88_ ( .D(Red_AddRoundKeyOutput[88]), 
        .CK(clk), .Q(Red_StateRegOutput[88]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_89_ ( .D(Red_AddRoundKeyOutput[89]), 
        .CK(clk), .Q(Red_StateRegOutput[89]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_90_ ( .D(Red_AddRoundKeyOutput[90]), 
        .CK(clk), .Q(Red_StateRegOutput[90]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_91_ ( .D(Red_AddRoundKeyOutput[91]), 
        .CK(clk), .Q(Red_StateRegOutput[91]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_92_ ( .D(Red_AddRoundKeyOutput[92]), 
        .CK(clk), .Q(Red_StateRegOutput[92]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_93_ ( .D(Red_AddRoundKeyOutput[93]), 
        .CK(clk), .Q(Red_StateRegOutput[93]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_94_ ( .D(Red_AddRoundKeyOutput[94]), 
        .CK(clk), .Q(Red_StateRegOutput[94]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_95_ ( .D(Red_AddRoundKeyOutput[95]), 
        .CK(clk), .Q(Red_StateRegOutput[95]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_96_ ( .D(Red_AddRoundKeyOutput[96]), 
        .CK(clk), .Q(Red_StateRegOutput[96]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_97_ ( .D(Red_AddRoundKeyOutput[97]), 
        .CK(clk), .Q(Red_StateRegOutput[97]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_98_ ( .D(Red_AddRoundKeyOutput[98]), 
        .CK(clk), .Q(Red_StateRegOutput[98]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_99_ ( .D(Red_AddRoundKeyOutput[99]), 
        .CK(clk), .Q(Red_StateRegOutput[99]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_100_ ( .D(Red_AddRoundKeyOutput[100]), .CK(clk), .Q(Red_StateRegOutput[100]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_101_ ( .D(Red_AddRoundKeyOutput[101]), .CK(clk), .Q(Red_StateRegOutput[101]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_102_ ( .D(Red_AddRoundKeyOutput[102]), .CK(clk), .Q(Red_StateRegOutput[102]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_103_ ( .D(Red_AddRoundKeyOutput[103]), .CK(clk), .Q(Red_StateRegOutput[103]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_104_ ( .D(Red_AddRoundKeyOutput[104]), .CK(clk), .Q(Red_StateRegOutput[104]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_105_ ( .D(Red_AddRoundKeyOutput[105]), .CK(clk), .Q(Red_StateRegOutput[105]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_106_ ( .D(Red_AddRoundKeyOutput[106]), .CK(clk), .Q(Red_StateRegOutput[106]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_107_ ( .D(Red_AddRoundKeyOutput[107]), .CK(clk), .Q(Red_StateRegOutput[107]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_108_ ( .D(Red_AddRoundKeyOutput[108]), .CK(clk), .Q(Red_StateRegOutput[108]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_109_ ( .D(Red_AddRoundKeyOutput[109]), .CK(clk), .Q(Red_StateRegOutput[109]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_110_ ( .D(Red_AddRoundKeyOutput[110]), .CK(clk), .Q(Red_StateRegOutput[110]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_111_ ( .D(Red_AddRoundKeyOutput[111]), .CK(clk), .Q(Red_StateRegOutput[111]), .QN() );
  BUF_X2 F_SD2_RedSB_inst_U64 ( .A(StateRegOutput[27]), .Z(
        F_SD2_RedSB_inst_n44) );
  BUF_X2 F_SD2_RedSB_inst_U63 ( .A(StateRegOutput[23]), .Z(
        F_SD2_RedSB_inst_n40) );
  BUF_X2 F_SD2_RedSB_inst_U62 ( .A(StateRegOutput[7]), .Z(F_SD2_RedSB_inst_n24) );
  BUF_X2 F_SD2_RedSB_inst_U61 ( .A(StateRegOutput[11]), .Z(
        F_SD2_RedSB_inst_n28) );
  BUF_X2 F_SD2_RedSB_inst_U60 ( .A(StateRegOutput[15]), .Z(
        F_SD2_RedSB_inst_n32) );
  BUF_X2 F_SD2_RedSB_inst_U59 ( .A(StateRegOutput[3]), .Z(F_SD2_RedSB_inst_n20) );
  BUF_X2 F_SD2_RedSB_inst_U58 ( .A(StateRegOutput[19]), .Z(
        F_SD2_RedSB_inst_n36) );
  BUF_X2 F_SD2_RedSB_inst_U57 ( .A(StateRegOutput[31]), .Z(
        F_SD2_RedSB_inst_n48) );
  BUF_X2 F_SD2_RedSB_inst_U56 ( .A(StateRegOutput[63]), .Z(
        F_SD2_RedSB_inst_n80) );
  BUF_X2 F_SD2_RedSB_inst_U55 ( .A(StateRegOutput[51]), .Z(
        F_SD2_RedSB_inst_n68) );
  BUF_X2 F_SD2_RedSB_inst_U54 ( .A(StateRegOutput[55]), .Z(
        F_SD2_RedSB_inst_n72) );
  BUF_X2 F_SD2_RedSB_inst_U53 ( .A(StateRegOutput[59]), .Z(
        F_SD2_RedSB_inst_n76) );
  BUF_X2 F_SD2_RedSB_inst_U52 ( .A(StateRegOutput[35]), .Z(
        F_SD2_RedSB_inst_n52) );
  BUF_X2 F_SD2_RedSB_inst_U51 ( .A(StateRegOutput[47]), .Z(
        F_SD2_RedSB_inst_n64) );
  BUF_X2 F_SD2_RedSB_inst_U50 ( .A(StateRegOutput[43]), .Z(
        F_SD2_RedSB_inst_n60) );
  BUF_X2 F_SD2_RedSB_inst_U49 ( .A(StateRegOutput[39]), .Z(
        F_SD2_RedSB_inst_n56) );
  BUF_X2 F_SD2_RedSB_inst_U48 ( .A(StateRegOutput[22]), .Z(
        F_SD2_RedSB_inst_n39) );
  BUF_X2 F_SD2_RedSB_inst_U47 ( .A(StateRegOutput[58]), .Z(
        F_SD2_RedSB_inst_n75) );
  BUF_X2 F_SD2_RedSB_inst_U46 ( .A(StateRegOutput[26]), .Z(
        F_SD2_RedSB_inst_n43) );
  BUF_X2 F_SD2_RedSB_inst_U45 ( .A(StateRegOutput[54]), .Z(
        F_SD2_RedSB_inst_n71) );
  BUF_X2 F_SD2_RedSB_inst_U44 ( .A(StateRegOutput[2]), .Z(F_SD2_RedSB_inst_n19) );
  BUF_X2 F_SD2_RedSB_inst_U43 ( .A(StateRegOutput[38]), .Z(
        F_SD2_RedSB_inst_n55) );
  BUF_X2 F_SD2_RedSB_inst_U42 ( .A(StateRegOutput[14]), .Z(
        F_SD2_RedSB_inst_n31) );
  BUF_X2 F_SD2_RedSB_inst_U41 ( .A(StateRegOutput[42]), .Z(
        F_SD2_RedSB_inst_n59) );
  BUF_X2 F_SD2_RedSB_inst_U40 ( .A(StateRegOutput[50]), .Z(
        F_SD2_RedSB_inst_n67) );
  BUF_X2 F_SD2_RedSB_inst_U39 ( .A(StateRegOutput[10]), .Z(
        F_SD2_RedSB_inst_n27) );
  BUF_X2 F_SD2_RedSB_inst_U38 ( .A(StateRegOutput[46]), .Z(
        F_SD2_RedSB_inst_n63) );
  BUF_X2 F_SD2_RedSB_inst_U37 ( .A(StateRegOutput[62]), .Z(
        F_SD2_RedSB_inst_n79) );
  BUF_X2 F_SD2_RedSB_inst_U36 ( .A(StateRegOutput[6]), .Z(F_SD2_RedSB_inst_n23) );
  BUF_X2 F_SD2_RedSB_inst_U35 ( .A(StateRegOutput[34]), .Z(
        F_SD2_RedSB_inst_n51) );
  BUF_X2 F_SD2_RedSB_inst_U34 ( .A(StateRegOutput[18]), .Z(
        F_SD2_RedSB_inst_n35) );
  BUF_X2 F_SD2_RedSB_inst_U33 ( .A(StateRegOutput[30]), .Z(
        F_SD2_RedSB_inst_n47) );
  BUF_X2 F_SD2_RedSB_inst_U32 ( .A(StateRegOutput[21]), .Z(
        F_SD2_RedSB_inst_n38) );
  BUF_X2 F_SD2_RedSB_inst_U31 ( .A(StateRegOutput[57]), .Z(
        F_SD2_RedSB_inst_n74) );
  BUF_X2 F_SD2_RedSB_inst_U30 ( .A(StateRegOutput[25]), .Z(
        F_SD2_RedSB_inst_n42) );
  BUF_X2 F_SD2_RedSB_inst_U29 ( .A(StateRegOutput[53]), .Z(
        F_SD2_RedSB_inst_n70) );
  BUF_X2 F_SD2_RedSB_inst_U28 ( .A(StateRegOutput[1]), .Z(F_SD2_RedSB_inst_n18) );
  BUF_X2 F_SD2_RedSB_inst_U27 ( .A(StateRegOutput[37]), .Z(
        F_SD2_RedSB_inst_n54) );
  BUF_X2 F_SD2_RedSB_inst_U26 ( .A(StateRegOutput[13]), .Z(
        F_SD2_RedSB_inst_n30) );
  BUF_X2 F_SD2_RedSB_inst_U25 ( .A(StateRegOutput[41]), .Z(
        F_SD2_RedSB_inst_n58) );
  BUF_X2 F_SD2_RedSB_inst_U24 ( .A(StateRegOutput[49]), .Z(
        F_SD2_RedSB_inst_n66) );
  BUF_X2 F_SD2_RedSB_inst_U23 ( .A(StateRegOutput[9]), .Z(F_SD2_RedSB_inst_n26) );
  BUF_X2 F_SD2_RedSB_inst_U22 ( .A(StateRegOutput[45]), .Z(
        F_SD2_RedSB_inst_n62) );
  BUF_X2 F_SD2_RedSB_inst_U21 ( .A(StateRegOutput[61]), .Z(
        F_SD2_RedSB_inst_n78) );
  BUF_X2 F_SD2_RedSB_inst_U20 ( .A(StateRegOutput[5]), .Z(F_SD2_RedSB_inst_n22) );
  BUF_X2 F_SD2_RedSB_inst_U19 ( .A(StateRegOutput[33]), .Z(
        F_SD2_RedSB_inst_n50) );
  BUF_X2 F_SD2_RedSB_inst_U18 ( .A(StateRegOutput[17]), .Z(
        F_SD2_RedSB_inst_n34) );
  BUF_X2 F_SD2_RedSB_inst_U17 ( .A(StateRegOutput[29]), .Z(
        F_SD2_RedSB_inst_n46) );
  BUF_X2 F_SD2_RedSB_inst_U16 ( .A(StateRegOutput[20]), .Z(
        F_SD2_RedSB_inst_n37) );
  BUF_X2 F_SD2_RedSB_inst_U15 ( .A(StateRegOutput[56]), .Z(
        F_SD2_RedSB_inst_n73) );
  BUF_X2 F_SD2_RedSB_inst_U14 ( .A(StateRegOutput[24]), .Z(
        F_SD2_RedSB_inst_n41) );
  BUF_X2 F_SD2_RedSB_inst_U13 ( .A(StateRegOutput[52]), .Z(
        F_SD2_RedSB_inst_n69) );
  BUF_X2 F_SD2_RedSB_inst_U12 ( .A(StateRegOutput[0]), .Z(F_SD2_RedSB_inst_n17) );
  BUF_X2 F_SD2_RedSB_inst_U11 ( .A(StateRegOutput[36]), .Z(
        F_SD2_RedSB_inst_n53) );
  BUF_X2 F_SD2_RedSB_inst_U10 ( .A(StateRegOutput[12]), .Z(
        F_SD2_RedSB_inst_n29) );
  BUF_X2 F_SD2_RedSB_inst_U9 ( .A(StateRegOutput[40]), .Z(F_SD2_RedSB_inst_n57) );
  BUF_X2 F_SD2_RedSB_inst_U8 ( .A(StateRegOutput[48]), .Z(F_SD2_RedSB_inst_n65) );
  BUF_X2 F_SD2_RedSB_inst_U7 ( .A(StateRegOutput[8]), .Z(F_SD2_RedSB_inst_n25)
         );
  BUF_X2 F_SD2_RedSB_inst_U6 ( .A(StateRegOutput[44]), .Z(F_SD2_RedSB_inst_n61) );
  BUF_X2 F_SD2_RedSB_inst_U5 ( .A(StateRegOutput[60]), .Z(F_SD2_RedSB_inst_n77) );
  BUF_X2 F_SD2_RedSB_inst_U4 ( .A(StateRegOutput[4]), .Z(F_SD2_RedSB_inst_n21)
         );
  BUF_X2 F_SD2_RedSB_inst_U3 ( .A(StateRegOutput[32]), .Z(F_SD2_RedSB_inst_n49) );
  BUF_X2 F_SD2_RedSB_inst_U2 ( .A(StateRegOutput[16]), .Z(F_SD2_RedSB_inst_n33) );
  BUF_X2 F_SD2_RedSB_inst_U1 ( .A(StateRegOutput[28]), .Z(F_SD2_RedSB_inst_n45) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_U69 ( .A(
        Red_StateRegOutput[1]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n280), .Z(Red_Feedback[105])
         );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_U68 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n279), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n278), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n280) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_U67 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n277), .B2(
        Red_StateRegOutput[2]), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n276), .C2(
        Red_StateRegOutput[5]), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n275), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n278) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_U66 ( .A1(
        Red_StateRegOutput[2]), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n277), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n276), .B2(
        Red_StateRegOutput[5]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n275) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_U65 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n274), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n273), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n276) );
  AOI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_U64 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n272), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n271), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n270), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n269), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n273) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_U63 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n268), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n267), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n266), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n265), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n264), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n269) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_U62 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n268), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n263), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n262), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n270) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_U61 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n268), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n263), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n261), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n262) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_U60 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n260), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n259), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n258), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n271) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_U59 ( .A(
        Red_StateRegOutput[0]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n257), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n274) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_U58 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n244), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n243), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n245), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n242), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n241), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n277) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_U57 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n240), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n239), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n238), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n241) );
  AOI222_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_U56 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n255), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n253), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n255), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n237), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n253), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n237), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n239) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_U55 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n247), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n267), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n237) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_U54 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n263), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n251), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n253) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_U53 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n236), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n255) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_U52 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n256), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n235), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n242) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_U51 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n261), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n263), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n234), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n243) );
  NOR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_U50 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n267), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n249), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n259), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n234) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_U49 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n250), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n251), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n259) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_U48 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n268), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n233), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n249) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_U47 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n256), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n267) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_U46 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n247), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n250), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n261) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_U45 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n264), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n260), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n232), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n279) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_U44 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n251), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n231), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n230), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n232) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_U43 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n251), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n229), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n252), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n230) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_U42 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n240), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n252) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_U41 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n247), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n265), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n240) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_U40 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n244), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n233), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n265) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_U39 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n246), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n248), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n256), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n263), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n229) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_U38 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n245), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n250), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n248) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_U37 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n266), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n247), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n246) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_U36 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n272), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n228), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n258), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n231) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_U35 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n236), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n227), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n258) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_U34 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n245), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n233), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n228) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_U33 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n236), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n227), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n260) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_U32 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n233), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n256), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n227) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_U31 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n226), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n225), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n256) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_U30 ( .A(
        Red_StateRegOutput[0]), .B(F_SD2_RedSB_inst_n17), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n226) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_U29 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n263), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n233) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_U28 ( .A(
        Red_StateRegOutput[6]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n224), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n263) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_U27 ( .A(
        F_SD2_RedSB_inst_n20), .B(F_SD2_RedSB_inst_n19), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n224) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_U26 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n244), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n268), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n236) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_U25 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n266), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n268) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_U24 ( .A(
        Red_StateRegOutput[4]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n225), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n266) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_U23 ( .A(
        F_SD2_RedSB_inst_n18), .B(F_SD2_RedSB_inst_n19), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n225) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_U22 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n245), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n244) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_U21 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n223), .B(
        Red_StateRegOutput[3]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n245) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_U20 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n235), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n264) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_U19 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n254), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n251), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n235) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_U18 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n222), .B(F_SD2_RedSB_inst_n18), .Z(F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n251) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_U17 ( .A(
        Red_StateRegOutput[1]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n223), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n222) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_U16 ( .A(
        F_SD2_RedSB_inst_n20), .B(F_SD2_RedSB_inst_n17), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n223) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_U15 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n247), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n250), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n254) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_U14 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n238), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n250) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_U13 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n221), .B(
        Red_StateRegOutput[2]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n238) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_U12 ( .A(
        F_SD2_RedSB_inst_n17), .B(F_SD2_RedSB_inst_n19), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n221) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_U11 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n272), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n247) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_U10 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n220), .B(F_SD2_RedSB_inst_n18), .ZN(F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n272) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_U9 ( .A(
        Red_StateRegOutput[5]), .B(F_SD2_RedSB_inst_n20), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n220) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_U8 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n215), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n217), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n256), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n219), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n257) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_U7 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n251), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n218), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n250), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n249), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n219) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_U6 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n247), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n248), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n245), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n246), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n218) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_U5 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n254), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n255), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n252), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n216), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n217) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_U4 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n267), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n216) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_U3 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n255), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n254), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n253), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_0_n215) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_U68 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n273), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n274) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_U67 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n272), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n271), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n275) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_U66 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n267), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n266), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n269) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_U65 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n272), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n271), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n264), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n265) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_U64 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n260), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n259), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n267), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n268), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n261) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_U63 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n258), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n257), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n268) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_U62 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n256), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n267), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n255), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n254), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n260) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_U61 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n253), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n267) );
  NOR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_U60 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n252), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n251), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n250), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n262) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_U59 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n270), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n263) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_U58 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n258), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n257), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n270) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_U57 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n272), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n249), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n257) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_U56 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n252), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n273), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n246) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_U55 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n264), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n250), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n273) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_U54 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n253), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n259), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n250) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_U53 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n266), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n264) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_U52 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n252), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n259), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n248) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_U51 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n278), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n259) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_U50 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n278), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n249), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n245) );
  AND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_U49 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n277), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n271), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n258) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_U48 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n272), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n253), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n255) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_U47 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n251), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n272) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_U46 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n251), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n277), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n256) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_U45 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n252), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n277) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_U44 ( .A(
        Red_StateRegOutput[5]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n244), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n278) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_U43 ( .A(
        F_SD2_RedSB_inst_n19), .B(F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n243), .ZN(F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n266) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_U42 ( .A(
        Red_StateRegOutput[2]), .B(F_SD2_RedSB_inst_n17), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n243) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_U41 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n254), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n276) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_U40 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n271), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n247), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n254) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_U39 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n249), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n247) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_U38 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n242), .B(
        Red_StateRegOutput[0]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n249) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_U37 ( .A(
        F_SD2_RedSB_inst_n17), .B(F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n241), .ZN(F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n242) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_U36 ( .A(
        Red_StateRegOutput[4]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n241), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n271) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_U35 ( .A(
        F_SD2_RedSB_inst_n19), .B(F_SD2_RedSB_inst_n18), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n241) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_U34 ( .A(
        Red_StateRegOutput[6]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n240), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n251) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_U33 ( .A(
        F_SD2_RedSB_inst_n19), .B(F_SD2_RedSB_inst_n20), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n240) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_U32 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n239), .B(
        Red_StateRegOutput[3]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n252) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_U31 ( .A(
        F_SD2_RedSB_inst_n17), .B(F_SD2_RedSB_inst_n20), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n239) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_U30 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n238), .B(
        Red_StateRegOutput[1]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n253) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_U29 ( .A(
        F_SD2_RedSB_inst_n17), .B(F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n244), .Z(F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n238) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_U28 ( .A(
        F_SD2_RedSB_inst_n18), .B(F_SD2_RedSB_inst_n20), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n244) );
  AOI222_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_U27 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n221), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n228), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n221), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n233), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n228), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n237), .ZN(Red_Feedback[106])
         );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_U26 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n236), .B(
        Red_StateRegOutput[1]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n237) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_U25 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n235), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n234), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n236) );
  NAND4_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_U24 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n249), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n252), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n264), .A4(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n255), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n235) );
  AOI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_U23 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n273), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n263), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n261), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n262), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n234) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_U22 ( .A(
        Red_StateRegOutput[5]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n232), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n233) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_U21 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n229), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n278), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n230), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n278), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n231), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n232) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_U20 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n277), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n276), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n275), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n276), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n274), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n231) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_U19 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n270), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n269), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n268), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n230) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_U18 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n272), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n271), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n265), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n229) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_U17 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n227), .B(
        Red_StateRegOutput[2]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n228) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_U16 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n266), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n222), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n226), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n227) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_U15 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n247), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n246), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n225), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n226) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_U14 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n224), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n255), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n224), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n245), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n264), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n225) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_U13 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n215), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n223), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n224) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_U12 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n251), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n248), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n258), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n245), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n223) );
  NOR4_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_U11 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n251), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n252), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n253), .A4(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n276), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n222) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_U10 ( .A(
        Red_StateRegOutput[0]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n220), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n221) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_U9 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n249), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n218), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n219), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n220) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_U8 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n249), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n215), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n214), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n219) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_U7 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n250), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n216), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n271), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n217), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n218) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_U6 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n264), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n272), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n253), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n248), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n217) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_U5 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n252), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n264), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n216) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_U4 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n278), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n256), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n258), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n255), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n215) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_U3 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n258), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n255), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n259), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n266), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_1_n214) );
  MUX2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_U54 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n240), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n239), .S(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n238), .Z(Red_Feedback[107])
         );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_U53 ( .A(
        Red_StateRegOutput[2]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n237), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n238) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_U52 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n236), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n235), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n234), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n233), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n237) );
  OR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_U51 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n232), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n231), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n230), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n233) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_U50 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n229), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n228), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n227), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n234) );
  AOI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_U49 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n226), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n225), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n224), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n223), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n236) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_U48 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n222), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n221), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n220), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n221), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n219), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n223) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_U47 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n226), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n225), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n218), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n221) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_U46 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n217), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n216), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n225) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_U45 ( .A(
        Red_StateRegOutput[5]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n215), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n239) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_U44 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n214), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n230), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n213), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n212), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n215) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_U43 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n228), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n226), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n211), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n232), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n212) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_U42 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n210), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n228), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n210), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n226), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n216), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n213) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_U41 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n220), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n216) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_U40 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n209), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n226) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_U39 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n208), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n207), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n228) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_U38 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n219), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n206), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n205), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n210) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_U37 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n219), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n206), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n208), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n205) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_U36 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n235), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n208) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_U35 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n222), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n204), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n229), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n214) );
  AND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_U34 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n206), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n219), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n204) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_U33 ( .A(
        Red_StateRegOutput[1]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n203), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n240) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_U32 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n202), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n201), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n200), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n201), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n199), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n203) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_U31 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n198), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n197), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n230), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n209), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n199) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_U30 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n227), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n220), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n218), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n197) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_U29 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n207), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n218) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_U28 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n222), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n201), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n227) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_U27 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n198), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n230), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n209), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n230), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n217), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n200) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_U26 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n231), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n206), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n209) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_U25 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n207), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n235), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n220), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n230) );
  AOI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_U24 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n229), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n211), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n207), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n224), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n198) );
  NOR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_U23 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n231), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n220), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n201), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n224) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_U22 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n219), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n220), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n211) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_U21 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n196), .B(
        Red_StateRegOutput[5]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n220) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_U20 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n201), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n219) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_U19 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n232), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n206), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n229) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_U18 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n195), .B(
        Red_StateRegOutput[4]), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n206) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_U17 ( .A(
        F_SD2_RedSB_inst_n19), .B(F_SD2_RedSB_inst_n18), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n195) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_U16 ( .A(
        Red_StateRegOutput[6]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n194), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n201) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_U15 ( .A(
        F_SD2_RedSB_inst_n19), .B(F_SD2_RedSB_inst_n20), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n194) );
  NOR4_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_U14 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n207), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n231), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n232), .A4(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n235), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n202) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_U13 ( .A(
        Red_StateRegOutput[2]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n193), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n235) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_U12 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n217), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n232) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_U11 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n192), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n193), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n217) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_U10 ( .A(
        F_SD2_RedSB_inst_n17), .B(F_SD2_RedSB_inst_n19), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n193) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_U9 ( .A(
        F_SD2_RedSB_inst_n18), .B(Red_StateRegOutput[0]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n192) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_U8 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n222), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n231) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_U7 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n191), .B(
        Red_StateRegOutput[3]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n222) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_U6 ( .A(
        F_SD2_RedSB_inst_n17), .B(F_SD2_RedSB_inst_n20), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n191) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_U5 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n190), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n196), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n207) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_U4 ( .A(F_SD2_RedSB_inst_n18), .B(F_SD2_RedSB_inst_n20), .Z(F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n196)
         );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_U3 ( .A(
        F_SD2_RedSB_inst_n17), .B(Red_StateRegOutput[1]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_2_n190) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_U70 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n290), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n289), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n288), .ZN(Red_Feedback[108])
         );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_U69 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n290), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n287), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n288) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_U68 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n286), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n285), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n284), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n287) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_U67 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n283), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n282), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n286), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n284) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_U66 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n289), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n285) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_U65 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n283), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n282), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n281), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n289) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_U64 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n282), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n286), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n283), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n281) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_U63 ( .A(
        Red_StateRegOutput[5]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n268), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n282) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_U62 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n267), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n266), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n265), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n269), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n268) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_U61 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n264), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n274), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n263), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n262), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n261), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n265) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_U60 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n260), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n259), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n278), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n258), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n263) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_U59 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n262), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n274) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_U58 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n273), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n272), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n264) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_U57 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n257), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n266) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_U56 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n256), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n255), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n254), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n267) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_U55 ( .A(
        Red_StateRegOutput[2]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n253), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n283) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_U54 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n252), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n262), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n251), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n250), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n253) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_U53 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n278), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n257), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n249), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n250) );
  NAND4_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_U52 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n254), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n248), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n276), .A4(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n262), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n251) );
  AOI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_U51 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n271), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n247), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n246), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n277), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n252) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_U50 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n258), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n259), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n245), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n277) );
  NOR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_U49 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n278), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n244), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n280), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n246) );
  AND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_U48 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n258), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n259), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n280) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_U47 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n243), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n259) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_U46 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n249), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n269), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n271) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_U45 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n276), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n279), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n257) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_U44 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n262), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n269), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n279) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_U43 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n244), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n256), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n245) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_U42 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n241), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n247), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n256) );
  AND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_U41 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n243), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n242), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n261) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_U40 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n278), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n272), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n242) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_U39 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n249), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n273), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n243) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_U38 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n255), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n273) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_U37 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n249), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n247), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n248) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_U36 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n275), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n255), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n254) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_U35 ( .A(
        Red_StateRegOutput[4]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n240), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n255) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_U34 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n278), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n275) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_U33 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n269), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n244) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_U32 ( .A(
        Red_StateRegOutput[5]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n239), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n269) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_U31 ( .A(
        F_SD2_RedSB_inst_n18), .B(F_SD2_RedSB_inst_n20), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n239) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_U30 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n262), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n241), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n270) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_U29 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n249), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n241) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_U28 ( .A(
        Red_StateRegOutput[3]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n238), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n249) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_U27 ( .A(
        F_SD2_RedSB_inst_n17), .B(F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n237), .ZN(F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n262) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_U26 ( .A(
        Red_StateRegOutput[2]), .B(F_SD2_RedSB_inst_n19), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n237) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_U25 ( .A(
        F_SD2_RedSB_inst_n18), .B(F_SD2_RedSB_inst_n19), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n240) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_U24 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n276), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n247), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n258) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_U23 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n272), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n247) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_U22 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n236), .B(
        Red_StateRegOutput[6]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n272) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_U21 ( .A(
        F_SD2_RedSB_inst_n19), .B(F_SD2_RedSB_inst_n20), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n236) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_U20 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n260), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n276) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_U19 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n235), .B(
        Red_StateRegOutput[1]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n260) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_U18 ( .A(
        F_SD2_RedSB_inst_n18), .B(F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n238), .Z(F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n235) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_U17 ( .A(
        F_SD2_RedSB_inst_n17), .B(F_SD2_RedSB_inst_n20), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n238) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_U16 ( .A(
        Red_StateRegOutput[1]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n234), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n290) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_U15 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n258), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n230), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n232), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n233), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n234) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_U14 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n261), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n269), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n261), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n248), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n260), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n233) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_U13 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n243), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n257), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n242), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n257), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n231), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n232) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_U12 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n260), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n245), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n231) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_U11 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n278), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n270), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n244), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n254), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n230) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_U10 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n229), .B(
        Red_StateRegOutput[0]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n286) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_U9 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n225), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n277), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n228), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n229) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_U8 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n276), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n226), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n275), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n227), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n228) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_U7 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n274), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n272), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n273), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n227) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_U6 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n269), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n270), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n273), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n271), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n226) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_U5 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n280), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n279), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n278), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n225) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_U4 ( .A(
        Red_StateRegOutput[0]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n224), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n278) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_U3 ( .A(F_SD2_RedSB_inst_n17), .B(F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n240), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_3_n224) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_U73 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n277), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n276), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n279), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n278) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_U72 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n275), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n274), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n273), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n277) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_U71 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n272), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n279) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_U70 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n266), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n265), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n264), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n267) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_U69 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n265), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n269) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_U68 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n280), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n263) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_U67 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n261), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n260), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n280) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_U66 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n264), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n281), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n258), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n276) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_U65 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n283), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n275), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n259) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_U64 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n264), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n257), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n283) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_U63 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n261), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n262), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n255), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n285), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n256) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_U62 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n272), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n254), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n285) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_U61 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n270), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n253), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n282) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_U60 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n286), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n274) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_U59 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n257), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n252), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n286) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_U58 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n260), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n271), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n251), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n249) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_U57 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n273), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n248), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n247), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n250) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_U56 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n284), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n247) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_U55 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n270), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n253), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n284) );
  OR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_U54 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n275), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n254), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n253) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_U53 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n266), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n270) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_U52 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n255), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n275), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n248) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_U51 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n281), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n255) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_U50 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n272), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n245), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n244), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n246) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_U49 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n260), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n262), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n243), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n242), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n244) );
  OR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_U48 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n251), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n271), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n268), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n242) );
  OR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_U47 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n281), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n254), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n261), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n268) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_U46 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n257), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n251) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_U45 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n266), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n252), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n265), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n241), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n254), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n243) );
  AND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_U44 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n266), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n252), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n241) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_U43 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n275), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n257), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n265) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_U42 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n264), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n281), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n252) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_U41 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n261), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n264) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_U40 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n272), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n273), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n266) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_U39 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n273), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n254), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n262) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_U38 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n271), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n273) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_U37 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n275), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n281), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n260) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_U36 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n258), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n275) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_U35 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n258), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n240), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n261), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n240), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n254), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n245) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_U34 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n239), .B(
        Red_StateRegOutput[0]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n254) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_U33 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n238), .B(F_SD2_RedSB_inst_n18), .ZN(F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n239) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_U32 ( .A(
        Red_StateRegOutput[2]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n238), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n261) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_U31 ( .A(
        F_SD2_RedSB_inst_n19), .B(F_SD2_RedSB_inst_n17), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n238) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_U30 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n257), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n281), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n271), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n240) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_U29 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n237), .B(
        Red_StateRegOutput[3]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n271) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_U28 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n236), .B(F_SD2_RedSB_inst_n18), .ZN(F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n281) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_U27 ( .A(
        Red_StateRegOutput[5]), .B(F_SD2_RedSB_inst_n20), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n236) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_U26 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n235), .B(
        Red_StateRegOutput[1]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n257) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_U25 ( .A(
        F_SD2_RedSB_inst_n18), .B(F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n237), .ZN(F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n235) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_U24 ( .A(
        F_SD2_RedSB_inst_n17), .B(F_SD2_RedSB_inst_n20), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n237) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_U23 ( .A(
        Red_StateRegOutput[6]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n234), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n258) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_U22 ( .A(
        F_SD2_RedSB_inst_n19), .B(F_SD2_RedSB_inst_n20), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n234) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_U21 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n233), .B(
        Red_StateRegOutput[4]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n272) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_U20 ( .A(
        F_SD2_RedSB_inst_n19), .B(F_SD2_RedSB_inst_n18), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n233) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_U19 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n217), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n221), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n231), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n225), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n232), .ZN(Red_Feedback[109])
         );
  NOR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_U18 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n221), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n225), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n231), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n232) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_U17 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n229), .B2(
        Red_StateRegOutput[2]), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n230), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n231) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_U16 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n229), .B2(
        Red_StateRegOutput[2]), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n217), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n230) );
  AOI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_U15 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n271), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n226), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n227), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n228), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n229) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_U14 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n262), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n286), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n271), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n263), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n228) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_U13 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n270), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n269), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n267), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n268), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n227) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_U12 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n285), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n259), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n276), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n226) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_U11 ( .A(
        Red_StateRegOutput[5]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n224), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n225) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_U10 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n285), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n286), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n222), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n223), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n224) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_U9 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n279), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n280), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n278), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n223) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_U8 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n284), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n282), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n284), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n283), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n281), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n222) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_U7 ( .A(
        Red_StateRegOutput[1]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n220), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n221) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_U6 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n219), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n218), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n220) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_U5 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n251), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n250), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n249), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n219) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_U4 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n265), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n256), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n282), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n274), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n218) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_U3 ( .A(
        Red_StateRegOutput[0]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n246), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_4_n217) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_U73 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n284), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n283), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n282), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n281), .ZN(Red_Feedback[110])
         );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_U72 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n280), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n281), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n279), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n283) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_U71 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n280), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n281), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n282), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n279) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_U70 ( .A(
        Red_StateRegOutput[5]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n278), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n282) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_U69 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n277), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n276), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n278) );
  NAND4_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_U68 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n275), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n274), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n273), .A4(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n272), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n276) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_U67 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n271), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n270), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n269), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n268), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n277) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_U66 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n267), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n268) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_U65 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n274), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n266), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n265), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n264), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n270) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_U64 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n263), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n265) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_U63 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n262), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n272), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n261), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n260), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n266) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_U62 ( .A(
        Red_StateRegOutput[1]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n259), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n281) );
  NOR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_U61 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n258), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n257), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n256), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n259) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_U60 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n255), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n254), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n255), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n253), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n252), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n256) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_U59 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n273), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n263), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n252) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_U58 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n251), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n250), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n263) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_U57 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n275), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n262), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n253) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_U56 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n271), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n269), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n254) );
  AOI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_U55 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n275), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n249), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n248), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n247), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n257) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_U54 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n246), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n245), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n275), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n247) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_U53 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n271), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n244), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n249) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_U52 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n245), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n271) );
  NOR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_U51 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n251), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n244), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n250), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n258) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_U50 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n260), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n248), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n250) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_U49 ( .A(
        Red_StateRegOutput[0]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n243), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n280) );
  AOI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_U48 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n275), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n242), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n241), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n240), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n243) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_U47 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n251), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n239), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n255), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n238), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n240) );
  OR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_U46 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n251), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n239), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n260), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n238) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_U45 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n237), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n248), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n244), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n255) );
  NOR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_U44 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n237), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n236), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n272), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n241) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_U43 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n274), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n262), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n246), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n235), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n236) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_U42 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n234), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n260), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n233), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n242) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_U41 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n232), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n246), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n262), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n233) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_U40 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n231), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n234) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_U39 ( .A(
        Red_StateRegOutput[2]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n230), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n284) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_U38 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n262), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n229), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n228), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n230) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_U37 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n267), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n227), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n226), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n264), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n228) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_U36 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n244), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n225), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n264) );
  NAND4_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_U35 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n237), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n269), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n274), .A4(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n227), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n226) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_U34 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n272), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n269) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_U33 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n237), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n273), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n262), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n231), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n267) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_U32 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n245), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n248), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n231) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_U31 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n244), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n239), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n273) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_U30 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n245), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n225), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n239) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_U29 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n260), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n237) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_U28 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n274), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n224), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n223), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n251), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n229) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_U27 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n232), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n244), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n261), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n244), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n235), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n224) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_U26 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n275), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n245), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n235) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_U25 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n227), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n275) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_U24 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n251), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n261) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_U23 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n227), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n272), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n251) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_U22 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n222), .B(
        Red_StateRegOutput[4]), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n272) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_U21 ( .A(
        F_SD2_RedSB_inst_n18), .B(F_SD2_RedSB_inst_n19), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n222) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_U20 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n221), .B(
        Red_StateRegOutput[3]), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n227) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_U19 ( .A(
        F_SD2_RedSB_inst_n17), .B(F_SD2_RedSB_inst_n20), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n221) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_U18 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n246), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n244) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_U17 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n220), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n219), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n246) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_U16 ( .A(
        F_SD2_RedSB_inst_n20), .B(Red_StateRegOutput[1]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n220) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_U15 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n223), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n232) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_U14 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n260), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n245), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n223) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_U13 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n218), .B(
        Red_StateRegOutput[5]), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n245) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_U12 ( .A(
        F_SD2_RedSB_inst_n18), .B(F_SD2_RedSB_inst_n20), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n218) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_U11 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n217), .B(F_SD2_RedSB_inst_n19), .Z(F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n260) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_U10 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n219), .B(
        Red_StateRegOutput[0]), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n217) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_U9 ( .A(
        F_SD2_RedSB_inst_n17), .B(F_SD2_RedSB_inst_n18), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n219) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_U8 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n248), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n274) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_U7 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n216), .B(
        Red_StateRegOutput[6]), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n248) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_U6 ( .A(
        F_SD2_RedSB_inst_n19), .B(F_SD2_RedSB_inst_n20), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n216) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_U5 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n225), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n262) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_U4 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n215), .B(F_SD2_RedSB_inst_n19), .Z(F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n225) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_U3 ( .A(
        Red_StateRegOutput[2]), .B(F_SD2_RedSB_inst_n17), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_5_n215) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_U65 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n176), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n175), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n174), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n173), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n172), .ZN(Red_Feedback[111])
         );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_U64 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n176), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n175), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n174), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n172) );
  MUX2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_U63 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n176), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n175), .S(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n171), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n173) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_U62 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n170), .B(
        Red_StateRegOutput[2]), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n171) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_U61 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n169), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n168), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n167), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n170) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_U60 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n166), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n167) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_U59 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n165), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n164), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n163), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n162), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n161), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n166) );
  AND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_U58 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n160), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n159), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n158), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n162) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_U57 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n159), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n157), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n156), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n155), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n168) );
  AOI222_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_U56 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n154), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n153), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n154), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n152), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n153), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n152), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n156) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_U55 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n151), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n161), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n152) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_U54 ( .A(
        Red_StateRegOutput[0]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n150), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n174) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_U53 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n161), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n149), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n148), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n150) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_U52 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n161), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n147), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n155), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n148) );
  AOI222_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_U51 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n154), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n153), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n154), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n146), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n153), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n146), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n147) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_U50 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n169), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n151), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n146) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_U49 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n145), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n144), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n143), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n142), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n149) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_U48 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n169), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n159), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n141), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n140), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n145) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_U47 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n157), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n140) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_U46 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n165), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n151), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n157) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_U45 ( .A(
        Red_StateRegOutput[1]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n139), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n175) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_U44 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n141), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n155), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n138), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n137), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n139) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_U43 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n141), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n136), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n137) );
  AOI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_U42 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n164), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n135), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n134), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n133), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n138) );
  NOR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_U41 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n163), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n132), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n143), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n133) );
  AND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_U40 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n131), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n161), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n153), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n134) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_U39 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n141), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n159), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n153) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_U38 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n144), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n130), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n142), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n131) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_U37 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n169), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n163), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n142) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_U36 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n151), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n129), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n155) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_U35 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n130), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n151) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_U34 ( .A(
        Red_StateRegOutput[5]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n128), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n176) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_U33 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n127), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n130), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n126), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n130), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n125), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n128) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_U32 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n144), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n161), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n160), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n129), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n164), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n125) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_U31 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n143), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n169), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n164) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_U30 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n130), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n141), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n143) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_U29 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n132), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n165), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n129) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_U28 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n135), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n158), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n136), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n126) );
  AND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_U27 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n154), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n124), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n136) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_U26 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n169), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n141), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n158) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_U25 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n123), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n122), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n141) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_U24 ( .A(
        F_SD2_RedSB_inst_n17), .B(Red_StateRegOutput[1]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n123) );
  OR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_U23 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n154), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n124), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n135) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_U22 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n161), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n159), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n124) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_U21 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n121), .B(
        Red_StateRegOutput[0]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n161) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_U20 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n120), .B(F_SD2_RedSB_inst_n18), .ZN(F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n121) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_U19 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n160), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n163), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n154) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_U18 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n165), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n163) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_U17 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n119), .B(
        Red_StateRegOutput[3]), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n165) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_U16 ( .A(
        F_SD2_RedSB_inst_n17), .B(F_SD2_RedSB_inst_n20), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n119) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_U15 ( .A(
        Red_StateRegOutput[5]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n122), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n130) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_U14 ( .A(
        F_SD2_RedSB_inst_n20), .B(F_SD2_RedSB_inst_n18), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n122) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_U13 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n118), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n127) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_U12 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n160), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n132), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n117), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n118) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_U11 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n160), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n132), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n169), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n117) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_U10 ( .A(
        Red_StateRegOutput[2]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n120), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n169) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_U9 ( .A(F_SD2_RedSB_inst_n19), .B(F_SD2_RedSB_inst_n17), .Z(F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n120)
         );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_U8 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n159), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n132) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_U7 ( .A(
        Red_StateRegOutput[6]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n116), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n159) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_U6 ( .A(F_SD2_RedSB_inst_n19), .B(F_SD2_RedSB_inst_n20), .Z(F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n116)
         );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_U5 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n144), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n160) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_U4 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n115), .B(
        Red_StateRegOutput[4]), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n144) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_U3 ( .A(
        F_SD2_RedSB_inst_n19), .B(F_SD2_RedSB_inst_n18), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_6_n115) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_U69 ( .A(
        Red_StateRegOutput[8]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n280), .Z(Red_Feedback[84]) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_U68 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n279), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n278), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n280) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_U67 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n277), .B2(
        Red_StateRegOutput[9]), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n276), .C2(
        Red_StateRegOutput[12]), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n275), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n278) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_U66 ( .A1(
        Red_StateRegOutput[9]), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n277), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n276), .B2(
        Red_StateRegOutput[12]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n275) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_U65 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n274), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n273), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n276) );
  AOI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_U64 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n272), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n271), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n270), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n269), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n273) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_U63 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n268), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n267), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n266), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n265), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n264), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n269) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_U62 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n268), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n263), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n262), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n270) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_U61 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n268), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n263), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n261), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n262) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_U60 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n260), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n259), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n258), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n271) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_U59 ( .A(
        Red_StateRegOutput[7]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n257), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n274) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_U58 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n244), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n243), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n245), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n242), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n241), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n277) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_U57 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n240), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n239), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n238), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n241) );
  AOI222_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_U56 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n255), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n253), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n255), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n237), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n253), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n237), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n239) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_U55 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n247), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n267), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n237) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_U54 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n263), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n251), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n253) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_U53 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n236), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n255) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_U52 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n256), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n235), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n242) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_U51 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n261), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n263), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n234), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n243) );
  NOR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_U50 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n267), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n249), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n259), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n234) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_U49 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n250), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n251), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n259) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_U48 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n268), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n233), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n249) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_U47 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n256), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n267) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_U46 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n247), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n250), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n261) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_U45 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n264), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n260), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n232), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n279) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_U44 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n251), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n231), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n230), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n232) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_U43 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n251), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n229), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n252), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n230) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_U42 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n240), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n252) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_U41 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n247), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n265), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n240) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_U40 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n244), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n233), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n265) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_U39 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n246), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n248), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n256), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n263), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n229) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_U38 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n245), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n250), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n248) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_U37 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n266), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n247), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n246) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_U36 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n272), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n228), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n258), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n231) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_U35 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n236), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n227), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n258) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_U34 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n245), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n233), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n228) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_U33 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n236), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n227), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n260) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_U32 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n233), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n256), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n227) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_U31 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n226), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n225), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n256) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_U30 ( .A(
        Red_StateRegOutput[7]), .B(F_SD2_RedSB_inst_n21), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n226) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_U29 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n263), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n233) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_U28 ( .A(
        Red_StateRegOutput[13]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n224), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n263) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_U27 ( .A(
        F_SD2_RedSB_inst_n24), .B(F_SD2_RedSB_inst_n23), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n224) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_U26 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n244), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n268), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n236) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_U25 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n266), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n268) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_U24 ( .A(
        Red_StateRegOutput[11]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n225), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n266) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_U23 ( .A(
        F_SD2_RedSB_inst_n22), .B(F_SD2_RedSB_inst_n23), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n225) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_U22 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n245), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n244) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_U21 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n223), .B(
        Red_StateRegOutput[10]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n245) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_U20 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n235), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n264) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_U19 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n254), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n251), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n235) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_U18 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n222), .B(F_SD2_RedSB_inst_n22), .Z(F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n251) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_U17 ( .A(
        Red_StateRegOutput[8]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n223), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n222) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_U16 ( .A(
        F_SD2_RedSB_inst_n24), .B(F_SD2_RedSB_inst_n21), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n223) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_U15 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n247), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n250), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n254) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_U14 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n238), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n250) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_U13 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n221), .B(
        Red_StateRegOutput[9]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n238) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_U12 ( .A(
        F_SD2_RedSB_inst_n21), .B(F_SD2_RedSB_inst_n23), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n221) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_U11 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n272), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n247) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_U10 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n220), .B(F_SD2_RedSB_inst_n22), .ZN(F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n272) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_U9 ( .A(
        Red_StateRegOutput[12]), .B(F_SD2_RedSB_inst_n24), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n220) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_U8 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n215), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n217), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n256), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n219), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n257) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_U7 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n251), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n218), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n250), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n249), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n219) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_U6 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n247), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n248), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n245), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n246), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n218) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_U5 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n254), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n255), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n252), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n216), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n217) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_U4 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n267), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n216) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_U3 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n255), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n254), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n253), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_7_n215) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_U68 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n273), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n274) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_U67 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n272), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n271), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n275) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_U66 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n267), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n266), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n269) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_U65 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n272), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n271), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n264), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n265) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_U64 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n260), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n259), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n267), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n268), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n261) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_U63 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n258), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n257), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n268) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_U62 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n256), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n267), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n255), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n254), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n260) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_U61 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n253), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n267) );
  NOR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_U60 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n252), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n251), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n250), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n262) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_U59 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n270), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n263) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_U58 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n258), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n257), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n270) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_U57 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n272), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n249), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n257) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_U56 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n252), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n273), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n246) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_U55 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n264), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n250), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n273) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_U54 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n253), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n259), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n250) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_U53 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n266), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n264) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_U52 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n252), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n259), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n248) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_U51 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n278), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n259) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_U50 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n278), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n249), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n245) );
  AND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_U49 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n277), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n271), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n258) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_U48 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n272), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n253), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n255) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_U47 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n251), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n272) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_U46 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n251), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n277), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n256) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_U45 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n252), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n277) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_U44 ( .A(
        Red_StateRegOutput[12]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n244), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n278) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_U43 ( .A(
        F_SD2_RedSB_inst_n23), .B(F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n243), .ZN(F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n266) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_U42 ( .A(
        Red_StateRegOutput[9]), .B(F_SD2_RedSB_inst_n21), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n243) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_U41 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n254), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n276) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_U40 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n271), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n247), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n254) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_U39 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n249), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n247) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_U38 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n242), .B(
        Red_StateRegOutput[7]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n249) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_U37 ( .A(
        F_SD2_RedSB_inst_n21), .B(F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n241), .ZN(F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n242) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_U36 ( .A(
        Red_StateRegOutput[11]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n241), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n271) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_U35 ( .A(
        F_SD2_RedSB_inst_n23), .B(F_SD2_RedSB_inst_n22), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n241) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_U34 ( .A(
        Red_StateRegOutput[13]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n240), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n251) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_U33 ( .A(
        F_SD2_RedSB_inst_n23), .B(F_SD2_RedSB_inst_n24), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n240) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_U32 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n239), .B(
        Red_StateRegOutput[10]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n252) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_U31 ( .A(
        F_SD2_RedSB_inst_n21), .B(F_SD2_RedSB_inst_n24), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n239) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_U30 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n238), .B(
        Red_StateRegOutput[8]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n253) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_U29 ( .A(
        F_SD2_RedSB_inst_n21), .B(F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n244), .Z(F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n238) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_U28 ( .A(
        F_SD2_RedSB_inst_n22), .B(F_SD2_RedSB_inst_n24), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n244) );
  AOI222_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_U27 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n221), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n228), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n221), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n233), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n228), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n237), .ZN(Red_Feedback[85])
         );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_U26 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n236), .B(
        Red_StateRegOutput[8]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n237) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_U25 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n234), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n235), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n236) );
  AOI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_U24 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n273), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n263), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n261), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n262), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n235) );
  NAND4_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_U23 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n249), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n252), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n264), .A4(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n255), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n234) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_U22 ( .A(
        Red_StateRegOutput[12]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n232), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n233) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_U21 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n229), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n278), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n230), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n278), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n231), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n232) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_U20 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n277), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n276), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n275), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n276), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n274), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n231) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_U19 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n270), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n269), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n268), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n230) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_U18 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n272), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n271), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n265), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n229) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_U17 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n227), .B(
        Red_StateRegOutput[9]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n228) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_U16 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n266), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n222), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n226), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n227) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_U15 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n247), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n246), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n225), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n226) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_U14 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n224), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n255), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n224), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n245), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n264), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n225) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_U13 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n217), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n223), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n224) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_U12 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n251), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n248), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n258), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n245), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n223) );
  NOR4_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_U11 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n251), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n252), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n253), .A4(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n276), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n222) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_U10 ( .A(
        Red_StateRegOutput[7]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n220), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n221) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_U9 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n249), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n216), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n219), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n220) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_U8 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n249), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n217), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n218), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n219) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_U7 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n258), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n255), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n259), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n266), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n218) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_U6 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n278), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n256), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n258), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n255), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n217) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_U5 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n250), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n214), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n271), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n215), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n216) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_U4 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n264), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n272), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n253), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n248), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n215) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_U3 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n252), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n264), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_8_n214) );
  MUX2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_U54 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n240), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n239), .S(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n238), .Z(Red_Feedback[86]) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_U53 ( .A(
        Red_StateRegOutput[9]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n237), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n238) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_U52 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n236), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n235), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n234), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n233), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n237) );
  OR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_U51 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n232), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n231), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n230), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n233) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_U50 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n229), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n228), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n227), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n234) );
  AOI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_U49 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n226), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n225), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n224), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n223), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n236) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_U48 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n222), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n221), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n220), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n221), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n219), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n223) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_U47 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n226), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n225), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n218), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n221) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_U46 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n217), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n216), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n225) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_U45 ( .A(
        Red_StateRegOutput[12]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n215), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n239) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_U44 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n214), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n230), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n213), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n212), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n215) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_U43 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n228), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n226), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n211), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n232), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n212) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_U42 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n210), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n228), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n210), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n226), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n216), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n213) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_U41 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n220), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n216) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_U40 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n209), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n226) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_U39 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n208), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n207), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n228) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_U38 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n219), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n206), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n205), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n210) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_U37 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n219), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n206), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n208), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n205) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_U36 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n235), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n208) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_U35 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n222), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n204), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n229), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n214) );
  AND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_U34 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n206), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n219), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n204) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_U33 ( .A(
        Red_StateRegOutput[8]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n203), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n240) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_U32 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n202), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n201), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n200), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n201), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n199), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n203) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_U31 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n198), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n197), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n230), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n209), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n199) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_U30 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n227), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n220), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n218), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n197) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_U29 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n207), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n218) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_U28 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n222), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n201), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n227) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_U27 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n198), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n230), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n209), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n230), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n217), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n200) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_U26 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n231), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n206), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n209) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_U25 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n207), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n235), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n220), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n230) );
  AOI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_U24 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n229), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n211), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n207), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n224), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n198) );
  NOR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_U23 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n231), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n220), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n201), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n224) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_U22 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n219), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n220), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n211) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_U21 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n196), .B(
        Red_StateRegOutput[12]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n220) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_U20 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n201), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n219) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_U19 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n232), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n206), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n229) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_U18 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n195), .B(
        Red_StateRegOutput[11]), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n206) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_U17 ( .A(
        F_SD2_RedSB_inst_n23), .B(F_SD2_RedSB_inst_n22), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n195) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_U16 ( .A(
        Red_StateRegOutput[13]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n194), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n201) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_U15 ( .A(
        F_SD2_RedSB_inst_n23), .B(F_SD2_RedSB_inst_n24), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n194) );
  NOR4_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_U14 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n207), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n231), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n232), .A4(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n235), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n202) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_U13 ( .A(
        Red_StateRegOutput[9]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n193), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n235) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_U12 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n217), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n232) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_U11 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n192), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n193), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n217) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_U10 ( .A(
        F_SD2_RedSB_inst_n21), .B(F_SD2_RedSB_inst_n23), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n193) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_U9 ( .A(
        F_SD2_RedSB_inst_n22), .B(Red_StateRegOutput[7]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n192) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_U8 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n222), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n231) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_U7 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n191), .B(
        Red_StateRegOutput[10]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n222) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_U6 ( .A(
        F_SD2_RedSB_inst_n21), .B(F_SD2_RedSB_inst_n24), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n191) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_U5 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n190), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n196), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n207) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_U4 ( .A(F_SD2_RedSB_inst_n22), .B(F_SD2_RedSB_inst_n24), .Z(F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n196)
         );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_U3 ( .A(
        F_SD2_RedSB_inst_n21), .B(Red_StateRegOutput[8]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_9_n190) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_U70 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n290), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n289), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n288), .ZN(Red_Feedback[87])
         );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_U69 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n290), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n287), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n288) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_U68 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n286), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n285), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n284), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n287) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_U67 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n283), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n282), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n286), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n284) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_U66 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n289), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n285) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_U65 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n283), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n282), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n281), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n289) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_U64 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n282), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n286), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n283), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n281) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_U63 ( .A(
        Red_StateRegOutput[12]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n268), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n282) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_U62 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n267), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n266), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n265), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n269), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n268) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_U61 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n264), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n274), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n263), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n262), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n261), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n265) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_U60 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n260), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n259), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n278), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n258), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n263) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_U59 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n262), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n274) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_U58 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n273), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n272), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n264) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_U57 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n257), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n266) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_U56 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n256), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n255), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n254), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n267) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_U55 ( .A(
        Red_StateRegOutput[9]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n253), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n283) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_U54 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n252), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n262), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n251), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n250), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n253) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_U53 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n278), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n257), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n249), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n250) );
  NAND4_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_U52 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n254), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n248), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n276), .A4(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n262), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n251) );
  AOI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_U51 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n271), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n247), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n246), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n277), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n252) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_U50 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n258), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n259), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n245), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n277) );
  NOR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_U49 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n278), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n244), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n280), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n246) );
  AND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_U48 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n258), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n259), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n280) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_U47 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n243), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n259) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_U46 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n249), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n269), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n271) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_U45 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n276), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n279), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n257) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_U44 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n262), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n269), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n279) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_U43 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n244), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n256), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n245) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_U42 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n241), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n247), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n256) );
  AND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_U41 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n243), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n242), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n261) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_U40 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n278), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n272), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n242) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_U39 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n249), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n273), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n243) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_U38 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n255), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n273) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_U37 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n249), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n247), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n248) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_U36 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n275), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n255), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n254) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_U35 ( .A(
        Red_StateRegOutput[11]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n240), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n255) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_U34 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n278), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n275) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_U33 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n269), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n244) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_U32 ( .A(
        Red_StateRegOutput[12]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n239), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n269) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_U31 ( .A(
        F_SD2_RedSB_inst_n22), .B(F_SD2_RedSB_inst_n24), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n239) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_U30 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n262), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n241), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n270) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_U29 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n249), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n241) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_U28 ( .A(
        Red_StateRegOutput[10]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n238), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n249) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_U27 ( .A(
        F_SD2_RedSB_inst_n21), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n237), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n262) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_U26 ( .A(
        Red_StateRegOutput[9]), .B(F_SD2_RedSB_inst_n23), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n237) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_U25 ( .A(
        F_SD2_RedSB_inst_n22), .B(F_SD2_RedSB_inst_n23), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n240) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_U24 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n276), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n247), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n258) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_U23 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n272), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n247) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_U22 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n236), .B(
        Red_StateRegOutput[13]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n272) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_U21 ( .A(
        F_SD2_RedSB_inst_n23), .B(F_SD2_RedSB_inst_n24), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n236) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_U20 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n260), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n276) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_U19 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n235), .B(
        Red_StateRegOutput[8]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n260) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_U18 ( .A(
        F_SD2_RedSB_inst_n22), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n238), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n235) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_U17 ( .A(
        F_SD2_RedSB_inst_n21), .B(F_SD2_RedSB_inst_n24), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n238) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_U16 ( .A(
        Red_StateRegOutput[8]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n234), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n290) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_U15 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n258), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n230), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n232), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n233), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n234) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_U14 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n261), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n269), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n261), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n248), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n260), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n233) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_U13 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n243), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n257), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n242), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n257), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n231), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n232) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_U12 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n260), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n245), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n231) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_U11 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n278), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n270), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n244), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n254), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n230) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_U10 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n229), .B(
        Red_StateRegOutput[7]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n286) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_U9 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n225), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n277), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n228), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n229) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_U8 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n276), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n226), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n275), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n227), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n228) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_U7 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n274), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n272), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n273), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n227) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_U6 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n269), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n270), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n273), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n271), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n226) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_U5 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n280), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n279), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n278), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n225) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_U4 ( .A(
        Red_StateRegOutput[7]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n224), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n278) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_U3 ( .A(
        F_SD2_RedSB_inst_n21), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n240), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_10_n224) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_U73 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n277), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n276), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n279), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n278) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_U72 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n275), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n274), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n273), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n277) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_U71 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n272), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n279) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_U70 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n266), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n265), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n264), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n267) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_U69 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n265), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n269) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_U68 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n280), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n263) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_U67 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n261), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n260), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n280) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_U66 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n264), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n281), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n258), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n276) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_U65 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n283), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n275), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n259) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_U64 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n264), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n257), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n283) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_U63 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n261), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n262), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n255), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n285), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n256) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_U62 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n272), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n254), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n285) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_U61 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n270), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n253), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n282) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_U60 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n286), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n274) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_U59 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n257), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n252), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n286) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_U58 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n260), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n271), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n251), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n249) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_U57 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n273), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n248), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n247), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n250) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_U56 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n284), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n247) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_U55 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n270), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n253), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n284) );
  OR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_U54 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n275), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n254), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n253) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_U53 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n266), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n270) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_U52 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n255), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n275), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n248) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_U51 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n281), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n255) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_U50 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n272), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n245), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n244), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n246) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_U49 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n260), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n262), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n243), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n242), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n244) );
  OR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_U48 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n251), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n271), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n268), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n242) );
  OR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_U47 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n281), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n254), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n261), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n268) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_U46 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n257), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n251) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_U45 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n266), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n252), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n265), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n241), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n254), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n243) );
  AND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_U44 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n266), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n252), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n241) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_U43 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n275), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n257), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n265) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_U42 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n264), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n281), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n252) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_U41 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n261), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n264) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_U40 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n272), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n273), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n266) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_U39 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n273), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n254), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n262) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_U38 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n271), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n273) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_U37 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n275), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n281), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n260) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_U36 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n258), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n275) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_U35 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n258), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n240), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n261), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n240), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n254), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n245) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_U34 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n239), .B(
        Red_StateRegOutput[7]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n254) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_U33 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n238), .B(
        F_SD2_RedSB_inst_n22), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n239) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_U32 ( .A(
        Red_StateRegOutput[9]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n238), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n261) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_U31 ( .A(
        F_SD2_RedSB_inst_n23), .B(F_SD2_RedSB_inst_n21), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n238) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_U30 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n257), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n281), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n271), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n240) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_U29 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n237), .B(
        Red_StateRegOutput[10]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n271) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_U28 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n236), .B(
        F_SD2_RedSB_inst_n22), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n281) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_U27 ( .A(
        Red_StateRegOutput[12]), .B(F_SD2_RedSB_inst_n24), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n236) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_U26 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n235), .B(
        Red_StateRegOutput[8]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n257) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_U25 ( .A(
        F_SD2_RedSB_inst_n22), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n237), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n235) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_U24 ( .A(
        F_SD2_RedSB_inst_n21), .B(F_SD2_RedSB_inst_n24), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n237) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_U23 ( .A(
        Red_StateRegOutput[13]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n234), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n258) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_U22 ( .A(
        F_SD2_RedSB_inst_n23), .B(F_SD2_RedSB_inst_n24), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n234) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_U21 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n233), .B(
        Red_StateRegOutput[11]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n272) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_U20 ( .A(
        F_SD2_RedSB_inst_n23), .B(F_SD2_RedSB_inst_n22), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n233) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_U19 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n217), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n221), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n227), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n231), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n232), .ZN(Red_Feedback[88])
         );
  NOR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_U18 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n221), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n231), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n227), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n232) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_U17 ( .A(
        Red_StateRegOutput[12]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n230), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n231) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_U16 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n285), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n286), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n228), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n229), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n230) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_U15 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n279), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n280), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n278), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n229) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_U14 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n284), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n282), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n284), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n283), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n281), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n228) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_U13 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n225), .B2(
        Red_StateRegOutput[9]), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n226), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n227) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_U12 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n225), .B2(
        Red_StateRegOutput[9]), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n217), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n226) );
  AOI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_U11 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n271), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n222), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n223), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n224), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n225) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_U10 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n262), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n286), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n271), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n263), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n224) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_U9 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n270), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n269), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n267), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n268), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n223) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_U8 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n285), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n259), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n276), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n222) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_U7 ( .A(
        Red_StateRegOutput[8]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n220), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n221) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_U6 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n218), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n219), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n220) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_U5 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n265), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n256), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n282), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n274), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n219) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_U4 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n251), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n250), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n249), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n218) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_U3 ( .A(
        Red_StateRegOutput[7]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n246), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_11_n217) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_U73 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n284), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n283), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n282), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n281), .ZN(Red_Feedback[89])
         );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_U72 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n280), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n281), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n279), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n283) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_U71 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n280), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n281), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n282), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n279) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_U70 ( .A(
        Red_StateRegOutput[12]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n278), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n282) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_U69 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n277), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n276), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n278) );
  NAND4_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_U68 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n275), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n274), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n273), .A4(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n272), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n276) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_U67 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n271), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n270), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n269), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n268), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n277) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_U66 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n267), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n268) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_U65 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n274), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n266), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n265), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n264), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n270) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_U64 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n263), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n265) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_U63 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n262), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n272), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n261), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n260), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n266) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_U62 ( .A(
        Red_StateRegOutput[8]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n259), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n281) );
  NOR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_U61 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n258), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n257), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n256), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n259) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_U60 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n255), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n254), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n255), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n253), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n252), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n256) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_U59 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n273), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n263), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n252) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_U58 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n251), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n250), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n263) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_U57 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n275), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n262), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n253) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_U56 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n271), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n269), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n254) );
  AOI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_U55 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n275), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n249), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n248), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n247), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n257) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_U54 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n246), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n245), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n275), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n247) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_U53 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n271), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n244), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n249) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_U52 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n245), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n271) );
  NOR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_U51 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n251), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n244), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n250), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n258) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_U50 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n260), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n248), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n250) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_U49 ( .A(
        Red_StateRegOutput[7]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n243), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n280) );
  AOI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_U48 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n275), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n242), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n241), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n240), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n243) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_U47 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n251), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n239), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n255), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n238), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n240) );
  OR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_U46 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n251), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n239), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n260), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n238) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_U45 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n237), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n248), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n244), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n255) );
  NOR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_U44 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n237), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n236), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n272), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n241) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_U43 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n274), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n262), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n246), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n235), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n236) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_U42 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n234), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n260), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n233), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n242) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_U41 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n232), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n246), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n262), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n233) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_U40 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n231), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n234) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_U39 ( .A(
        Red_StateRegOutput[9]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n230), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n284) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_U38 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n262), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n229), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n228), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n230) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_U37 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n267), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n227), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n226), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n264), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n228) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_U36 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n244), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n225), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n264) );
  NAND4_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_U35 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n237), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n269), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n274), .A4(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n227), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n226) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_U34 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n272), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n269) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_U33 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n237), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n273), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n262), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n231), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n267) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_U32 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n245), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n248), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n231) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_U31 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n244), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n239), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n273) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_U30 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n245), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n225), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n239) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_U29 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n260), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n237) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_U28 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n274), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n224), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n223), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n251), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n229) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_U27 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n232), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n244), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n261), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n244), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n235), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n224) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_U26 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n275), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n245), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n235) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_U25 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n227), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n275) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_U24 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n251), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n261) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_U23 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n227), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n272), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n251) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_U22 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n222), .B(
        Red_StateRegOutput[11]), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n272) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_U21 ( .A(
        F_SD2_RedSB_inst_n22), .B(F_SD2_RedSB_inst_n23), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n222) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_U20 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n221), .B(
        Red_StateRegOutput[10]), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n227) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_U19 ( .A(
        F_SD2_RedSB_inst_n21), .B(F_SD2_RedSB_inst_n24), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n221) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_U18 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n246), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n244) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_U17 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n220), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n219), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n246) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_U16 ( .A(
        F_SD2_RedSB_inst_n24), .B(Red_StateRegOutput[8]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n220) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_U15 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n223), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n232) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_U14 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n260), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n245), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n223) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_U13 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n218), .B(
        Red_StateRegOutput[12]), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n245) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_U12 ( .A(
        F_SD2_RedSB_inst_n22), .B(F_SD2_RedSB_inst_n24), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n218) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_U11 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n217), .B(
        F_SD2_RedSB_inst_n23), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n260) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_U10 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n219), .B(
        Red_StateRegOutput[7]), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n217) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_U9 ( .A(
        F_SD2_RedSB_inst_n21), .B(F_SD2_RedSB_inst_n22), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n219) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_U8 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n248), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n274) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_U7 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n216), .B(
        Red_StateRegOutput[13]), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n248) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_U6 ( .A(
        F_SD2_RedSB_inst_n23), .B(F_SD2_RedSB_inst_n24), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n216) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_U5 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n225), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n262) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_U4 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n215), .B(
        F_SD2_RedSB_inst_n23), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n225) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_U3 ( .A(
        Red_StateRegOutput[9]), .B(F_SD2_RedSB_inst_n21), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_12_n215) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_U65 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n283), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n282), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n281), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n280), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n279), .ZN(Red_Feedback[90])
         );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_U64 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n283), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n282), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n281), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n279) );
  MUX2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_U63 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n283), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n282), .S(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n278), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n280) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_U62 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n277), .B(
        Red_StateRegOutput[9]), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n278) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_U61 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n276), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n275), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n274), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n277) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_U60 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n273), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n274) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_U59 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n272), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n271), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n270), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n269), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n268), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n273) );
  AND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_U58 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n267), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n266), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n265), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n269) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_U57 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n266), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n264), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n263), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n262), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n275) );
  AOI222_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_U56 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n261), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n260), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n261), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n259), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n260), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n259), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n263) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_U55 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n258), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n268), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n259) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_U54 ( .A(
        Red_StateRegOutput[7]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n257), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n281) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_U53 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n268), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n256), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n255), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n257) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_U52 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n268), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n254), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n262), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n255) );
  AOI222_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_U51 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n261), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n260), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n261), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n253), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n260), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n253), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n254) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_U50 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n276), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n258), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n253) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_U49 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n252), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n251), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n250), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n249), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n256) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_U48 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n276), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n266), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n248), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n247), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n252) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_U47 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n264), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n247) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_U46 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n272), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n258), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n264) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_U45 ( .A(
        Red_StateRegOutput[8]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n246), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n282) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_U44 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n248), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n262), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n245), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n244), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n246) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_U43 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n248), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n243), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n244) );
  AOI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_U42 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n271), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n242), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n241), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n240), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n245) );
  NOR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_U41 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n270), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n239), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n250), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n240) );
  AND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_U40 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n238), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n268), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n260), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n241) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_U39 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n248), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n266), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n260) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_U38 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n251), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n237), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n249), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n238) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_U37 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n276), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n270), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n249) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_U36 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n258), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n236), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n262) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_U35 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n237), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n258) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_U34 ( .A(
        Red_StateRegOutput[12]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n235), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n283) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_U33 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n234), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n237), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n233), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n237), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n232), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n235) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_U32 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n251), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n268), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n267), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n236), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n271), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n232) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_U31 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n250), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n276), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n271) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_U30 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n237), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n248), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n250) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_U29 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n239), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n272), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n236) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_U28 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n242), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n265), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n243), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n233) );
  AND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_U27 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n261), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n231), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n243) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_U26 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n276), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n248), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n265) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_U25 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n230), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n229), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n248) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_U24 ( .A(
        F_SD2_RedSB_inst_n21), .B(Red_StateRegOutput[8]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n230) );
  OR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_U23 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n261), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n231), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n242) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_U22 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n268), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n266), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n231) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_U21 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n228), .B(
        Red_StateRegOutput[7]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n268) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_U20 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n227), .B(
        F_SD2_RedSB_inst_n22), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n228) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_U19 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n267), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n270), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n261) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_U18 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n272), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n270) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_U17 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n226), .B(
        Red_StateRegOutput[10]), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n272) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_U16 ( .A(
        F_SD2_RedSB_inst_n21), .B(F_SD2_RedSB_inst_n24), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n226) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_U15 ( .A(
        Red_StateRegOutput[12]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n229), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n237) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_U14 ( .A(
        F_SD2_RedSB_inst_n24), .B(F_SD2_RedSB_inst_n22), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n229) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_U13 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n225), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n234) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_U12 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n267), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n239), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n224), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n225) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_U11 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n267), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n239), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n276), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n224) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_U10 ( .A(
        Red_StateRegOutput[9]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n227), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n276) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_U9 ( .A(
        F_SD2_RedSB_inst_n23), .B(F_SD2_RedSB_inst_n21), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n227) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_U8 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n266), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n239) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_U7 ( .A(
        Red_StateRegOutput[13]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n223), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n266) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_U6 ( .A(
        F_SD2_RedSB_inst_n23), .B(F_SD2_RedSB_inst_n24), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n223) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_U5 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n251), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n267) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_U4 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n222), .B(
        Red_StateRegOutput[11]), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n251) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_U3 ( .A(
        F_SD2_RedSB_inst_n23), .B(F_SD2_RedSB_inst_n22), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_13_n222) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_U69 ( .A(
        Red_StateRegOutput[15]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n280), .Z(Red_Feedback[91])
         );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_U68 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n279), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n278), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n280) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_U67 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n277), .B2(
        Red_StateRegOutput[16]), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n276), .C2(
        Red_StateRegOutput[19]), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n275), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n278) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_U66 ( .A1(
        Red_StateRegOutput[16]), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n277), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n276), .B2(
        Red_StateRegOutput[19]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n275) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_U65 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n274), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n273), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n276) );
  AOI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_U64 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n272), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n271), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n270), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n269), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n273) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_U63 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n268), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n267), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n266), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n265), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n264), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n269) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_U62 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n268), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n263), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n262), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n270) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_U61 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n268), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n263), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n261), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n262) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_U60 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n260), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n259), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n258), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n271) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_U59 ( .A(
        Red_StateRegOutput[14]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n257), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n274) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_U58 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n244), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n243), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n245), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n242), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n241), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n277) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_U57 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n240), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n239), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n238), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n241) );
  AOI222_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_U56 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n255), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n253), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n255), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n237), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n253), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n237), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n239) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_U55 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n247), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n267), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n237) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_U54 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n263), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n251), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n253) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_U53 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n236), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n255) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_U52 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n256), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n235), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n242) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_U51 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n261), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n263), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n234), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n243) );
  NOR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_U50 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n267), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n249), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n259), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n234) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_U49 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n250), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n251), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n259) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_U48 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n268), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n233), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n249) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_U47 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n256), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n267) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_U46 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n247), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n250), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n261) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_U45 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n264), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n260), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n232), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n279) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_U44 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n251), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n231), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n230), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n232) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_U43 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n251), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n229), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n252), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n230) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_U42 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n240), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n252) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_U41 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n247), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n265), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n240) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_U40 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n244), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n233), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n265) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_U39 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n246), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n248), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n256), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n263), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n229) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_U38 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n245), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n250), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n248) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_U37 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n266), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n247), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n246) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_U36 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n272), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n228), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n258), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n231) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_U35 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n236), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n227), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n258) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_U34 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n245), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n233), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n228) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_U33 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n236), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n227), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n260) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_U32 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n233), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n256), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n227) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_U31 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n226), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n225), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n256) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_U30 ( .A(
        Red_StateRegOutput[14]), .B(F_SD2_RedSB_inst_n25), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n226) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_U29 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n263), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n233) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_U28 ( .A(
        Red_StateRegOutput[20]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n224), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n263) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_U27 ( .A(
        F_SD2_RedSB_inst_n28), .B(F_SD2_RedSB_inst_n27), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n224) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_U26 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n244), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n268), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n236) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_U25 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n266), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n268) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_U24 ( .A(
        Red_StateRegOutput[18]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n225), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n266) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_U23 ( .A(
        F_SD2_RedSB_inst_n26), .B(F_SD2_RedSB_inst_n27), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n225) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_U22 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n245), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n244) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_U21 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n223), .B(
        Red_StateRegOutput[17]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n245) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_U20 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n235), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n264) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_U19 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n254), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n251), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n235) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_U18 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n222), .B(
        F_SD2_RedSB_inst_n26), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n251) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_U17 ( .A(
        Red_StateRegOutput[15]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n223), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n222) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_U16 ( .A(
        F_SD2_RedSB_inst_n28), .B(F_SD2_RedSB_inst_n25), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n223) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_U15 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n247), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n250), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n254) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_U14 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n238), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n250) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_U13 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n221), .B(
        Red_StateRegOutput[16]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n238) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_U12 ( .A(
        F_SD2_RedSB_inst_n25), .B(F_SD2_RedSB_inst_n27), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n221) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_U11 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n272), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n247) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_U10 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n220), .B(
        F_SD2_RedSB_inst_n26), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n272) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_U9 ( .A(
        Red_StateRegOutput[19]), .B(F_SD2_RedSB_inst_n28), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n220) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_U8 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n215), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n217), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n256), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n219), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n257) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_U7 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n251), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n218), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n250), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n249), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n219) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_U6 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n247), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n248), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n245), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n246), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n218) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_U5 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n254), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n255), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n252), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n216), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n217) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_U4 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n267), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n216) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_U3 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n255), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n254), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n253), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_14_n215) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_U68 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n273), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n274) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_U67 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n272), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n271), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n275) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_U66 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n267), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n266), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n269) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_U65 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n272), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n271), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n264), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n265) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_U64 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n260), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n259), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n267), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n268), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n261) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_U63 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n258), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n257), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n268) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_U62 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n256), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n267), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n255), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n254), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n260) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_U61 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n253), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n267) );
  NOR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_U60 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n252), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n251), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n250), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n262) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_U59 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n270), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n263) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_U58 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n258), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n257), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n270) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_U57 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n272), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n249), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n257) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_U56 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n252), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n273), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n246) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_U55 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n264), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n250), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n273) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_U54 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n253), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n259), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n250) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_U53 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n266), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n264) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_U52 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n252), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n259), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n248) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_U51 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n278), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n259) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_U50 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n278), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n249), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n245) );
  AND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_U49 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n277), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n271), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n258) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_U48 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n272), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n253), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n255) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_U47 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n251), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n272) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_U46 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n251), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n277), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n256) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_U45 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n252), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n277) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_U44 ( .A(
        Red_StateRegOutput[19]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n244), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n278) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_U43 ( .A(
        F_SD2_RedSB_inst_n27), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n243), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n266) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_U42 ( .A(
        Red_StateRegOutput[16]), .B(F_SD2_RedSB_inst_n25), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n243) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_U41 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n254), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n276) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_U40 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n271), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n247), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n254) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_U39 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n249), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n247) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_U38 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n242), .B(
        Red_StateRegOutput[14]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n249) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_U37 ( .A(
        F_SD2_RedSB_inst_n25), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n241), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n242) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_U36 ( .A(
        Red_StateRegOutput[18]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n241), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n271) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_U35 ( .A(
        F_SD2_RedSB_inst_n27), .B(F_SD2_RedSB_inst_n26), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n241) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_U34 ( .A(
        Red_StateRegOutput[20]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n240), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n251) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_U33 ( .A(
        F_SD2_RedSB_inst_n27), .B(F_SD2_RedSB_inst_n28), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n240) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_U32 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n239), .B(
        Red_StateRegOutput[17]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n252) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_U31 ( .A(
        F_SD2_RedSB_inst_n25), .B(F_SD2_RedSB_inst_n28), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n239) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_U30 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n238), .B(
        Red_StateRegOutput[15]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n253) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_U29 ( .A(
        F_SD2_RedSB_inst_n25), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n244), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n238) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_U28 ( .A(
        F_SD2_RedSB_inst_n26), .B(F_SD2_RedSB_inst_n28), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n244) );
  AOI222_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_U27 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n221), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n228), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n221), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n233), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n228), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n237), .ZN(Red_Feedback[92])
         );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_U26 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n236), .B(
        Red_StateRegOutput[15]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n237) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_U25 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n234), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n235), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n236) );
  AOI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_U24 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n273), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n263), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n261), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n262), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n235) );
  NAND4_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_U23 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n249), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n252), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n264), .A4(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n255), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n234) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_U22 ( .A(
        Red_StateRegOutput[19]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n232), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n233) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_U21 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n229), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n278), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n230), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n278), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n231), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n232) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_U20 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n277), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n276), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n275), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n276), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n274), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n231) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_U19 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n270), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n269), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n268), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n230) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_U18 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n272), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n271), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n265), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n229) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_U17 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n227), .B(
        Red_StateRegOutput[16]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n228) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_U16 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n266), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n222), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n226), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n227) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_U15 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n247), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n246), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n225), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n226) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_U14 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n224), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n255), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n224), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n245), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n264), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n225) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_U13 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n217), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n223), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n224) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_U12 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n251), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n248), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n258), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n245), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n223) );
  NOR4_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_U11 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n251), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n252), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n253), .A4(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n276), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n222) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_U10 ( .A(
        Red_StateRegOutput[14]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n220), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n221) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_U9 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n249), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n216), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n219), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n220) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_U8 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n249), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n217), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n218), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n219) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_U7 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n258), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n255), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n259), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n266), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n218) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_U6 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n278), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n256), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n258), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n255), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n217) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_U5 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n250), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n214), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n271), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n215), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n216) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_U4 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n264), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n272), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n253), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n248), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n215) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_U3 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n252), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n264), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_15_n214) );
  MUX2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_U54 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n240), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n239), .S(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n238), .Z(Red_Feedback[93])
         );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_U53 ( .A(
        Red_StateRegOutput[16]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n237), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n238) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_U52 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n236), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n235), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n234), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n233), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n237) );
  OR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_U51 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n232), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n231), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n230), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n233) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_U50 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n229), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n228), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n227), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n234) );
  AOI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_U49 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n226), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n225), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n224), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n223), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n236) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_U48 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n222), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n221), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n220), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n221), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n219), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n223) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_U47 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n226), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n225), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n218), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n221) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_U46 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n217), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n216), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n225) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_U45 ( .A(
        Red_StateRegOutput[19]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n215), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n239) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_U44 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n214), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n230), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n213), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n212), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n215) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_U43 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n228), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n226), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n211), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n232), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n212) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_U42 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n210), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n228), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n210), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n226), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n216), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n213) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_U41 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n220), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n216) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_U40 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n209), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n226) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_U39 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n208), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n207), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n228) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_U38 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n219), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n206), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n205), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n210) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_U37 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n219), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n206), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n208), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n205) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_U36 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n235), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n208) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_U35 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n222), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n204), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n229), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n214) );
  AND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_U34 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n206), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n219), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n204) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_U33 ( .A(
        Red_StateRegOutput[15]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n203), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n240) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_U32 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n202), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n201), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n200), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n201), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n199), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n203) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_U31 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n198), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n197), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n230), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n209), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n199) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_U30 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n227), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n220), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n218), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n197) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_U29 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n207), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n218) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_U28 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n222), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n201), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n227) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_U27 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n198), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n230), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n209), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n230), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n217), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n200) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_U26 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n231), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n206), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n209) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_U25 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n207), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n235), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n220), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n230) );
  AOI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_U24 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n229), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n211), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n207), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n224), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n198) );
  NOR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_U23 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n231), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n220), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n201), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n224) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_U22 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n219), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n220), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n211) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_U21 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n196), .B(
        Red_StateRegOutput[19]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n220) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_U20 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n201), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n219) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_U19 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n232), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n206), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n229) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_U18 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n195), .B(
        Red_StateRegOutput[18]), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n206) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_U17 ( .A(
        F_SD2_RedSB_inst_n27), .B(F_SD2_RedSB_inst_n26), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n195) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_U16 ( .A(
        Red_StateRegOutput[20]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n194), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n201) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_U15 ( .A(
        F_SD2_RedSB_inst_n27), .B(F_SD2_RedSB_inst_n28), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n194) );
  NOR4_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_U14 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n207), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n231), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n232), .A4(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n235), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n202) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_U13 ( .A(
        Red_StateRegOutput[16]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n193), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n235) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_U12 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n217), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n232) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_U11 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n192), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n193), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n217) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_U10 ( .A(
        F_SD2_RedSB_inst_n25), .B(F_SD2_RedSB_inst_n27), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n193) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_U9 ( .A(
        F_SD2_RedSB_inst_n26), .B(Red_StateRegOutput[14]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n192) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_U8 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n222), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n231) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_U7 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n191), .B(
        Red_StateRegOutput[17]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n222) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_U6 ( .A(
        F_SD2_RedSB_inst_n25), .B(F_SD2_RedSB_inst_n28), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n191) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_U5 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n190), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n196), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n207) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_U4 ( .A(
        F_SD2_RedSB_inst_n26), .B(F_SD2_RedSB_inst_n28), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n196) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_U3 ( .A(
        F_SD2_RedSB_inst_n25), .B(Red_StateRegOutput[15]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_16_n190) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_U70 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n290), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n289), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n288), .ZN(Red_Feedback[94])
         );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_U69 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n290), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n287), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n288) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_U68 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n286), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n285), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n284), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n287) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_U67 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n283), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n282), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n286), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n284) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_U66 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n289), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n285) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_U65 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n283), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n282), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n281), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n289) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_U64 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n282), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n286), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n283), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n281) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_U63 ( .A(
        Red_StateRegOutput[19]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n268), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n282) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_U62 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n267), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n266), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n265), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n269), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n268) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_U61 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n264), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n274), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n263), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n262), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n261), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n265) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_U60 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n260), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n259), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n278), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n258), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n263) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_U59 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n262), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n274) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_U58 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n273), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n272), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n264) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_U57 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n257), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n266) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_U56 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n256), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n255), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n254), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n267) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_U55 ( .A(
        Red_StateRegOutput[16]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n253), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n283) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_U54 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n252), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n262), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n251), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n250), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n253) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_U53 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n278), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n257), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n249), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n250) );
  NAND4_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_U52 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n254), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n248), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n276), .A4(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n262), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n251) );
  AOI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_U51 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n271), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n247), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n246), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n277), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n252) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_U50 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n258), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n259), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n245), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n277) );
  NOR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_U49 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n278), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n244), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n280), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n246) );
  AND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_U48 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n258), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n259), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n280) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_U47 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n243), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n259) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_U46 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n249), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n269), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n271) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_U45 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n276), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n279), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n257) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_U44 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n262), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n269), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n279) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_U43 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n244), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n256), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n245) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_U42 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n241), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n247), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n256) );
  AND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_U41 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n243), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n242), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n261) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_U40 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n278), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n272), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n242) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_U39 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n249), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n273), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n243) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_U38 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n255), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n273) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_U37 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n249), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n247), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n248) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_U36 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n275), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n255), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n254) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_U35 ( .A(
        Red_StateRegOutput[18]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n240), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n255) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_U34 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n278), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n275) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_U33 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n269), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n244) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_U32 ( .A(
        Red_StateRegOutput[19]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n239), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n269) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_U31 ( .A(
        F_SD2_RedSB_inst_n26), .B(F_SD2_RedSB_inst_n28), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n239) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_U30 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n262), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n241), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n270) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_U29 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n249), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n241) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_U28 ( .A(
        Red_StateRegOutput[17]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n238), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n249) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_U27 ( .A(
        F_SD2_RedSB_inst_n25), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n237), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n262) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_U26 ( .A(
        Red_StateRegOutput[16]), .B(F_SD2_RedSB_inst_n27), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n237) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_U25 ( .A(
        F_SD2_RedSB_inst_n26), .B(F_SD2_RedSB_inst_n27), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n240) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_U24 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n276), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n247), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n258) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_U23 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n272), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n247) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_U22 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n236), .B(
        Red_StateRegOutput[20]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n272) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_U21 ( .A(
        F_SD2_RedSB_inst_n27), .B(F_SD2_RedSB_inst_n28), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n236) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_U20 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n260), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n276) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_U19 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n235), .B(
        Red_StateRegOutput[15]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n260) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_U18 ( .A(
        F_SD2_RedSB_inst_n26), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n238), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n235) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_U17 ( .A(
        F_SD2_RedSB_inst_n25), .B(F_SD2_RedSB_inst_n28), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n238) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_U16 ( .A(
        Red_StateRegOutput[15]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n234), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n290) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_U15 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n258), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n230), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n232), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n233), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n234) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_U14 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n261), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n269), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n261), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n248), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n260), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n233) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_U13 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n243), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n257), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n242), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n257), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n231), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n232) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_U12 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n260), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n245), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n231) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_U11 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n278), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n270), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n244), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n254), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n230) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_U10 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n229), .B(
        Red_StateRegOutput[14]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n286) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_U9 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n225), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n277), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n228), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n229) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_U8 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n276), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n226), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n275), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n227), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n228) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_U7 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n274), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n272), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n273), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n227) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_U6 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n269), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n270), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n273), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n271), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n226) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_U5 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n280), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n279), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n278), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n225) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_U4 ( .A(
        Red_StateRegOutput[14]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n224), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n278) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_U3 ( .A(
        F_SD2_RedSB_inst_n25), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n240), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_17_n224) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_U73 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n277), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n276), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n279), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n278) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_U72 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n275), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n274), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n273), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n277) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_U71 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n272), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n279) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_U70 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n266), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n265), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n264), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n267) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_U69 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n265), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n269) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_U68 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n280), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n263) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_U67 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n261), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n260), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n280) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_U66 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n264), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n281), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n258), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n276) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_U65 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n283), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n275), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n259) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_U64 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n264), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n257), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n283) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_U63 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n261), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n262), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n255), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n285), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n256) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_U62 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n272), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n254), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n285) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_U61 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n270), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n253), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n282) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_U60 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n286), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n274) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_U59 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n257), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n252), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n286) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_U58 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n260), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n271), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n251), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n249) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_U57 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n273), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n248), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n247), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n250) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_U56 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n284), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n247) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_U55 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n270), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n253), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n284) );
  OR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_U54 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n275), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n254), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n253) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_U53 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n266), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n270) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_U52 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n255), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n275), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n248) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_U51 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n281), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n255) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_U50 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n272), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n245), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n244), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n246) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_U49 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n260), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n262), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n243), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n242), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n244) );
  OR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_U48 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n251), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n271), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n268), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n242) );
  OR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_U47 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n281), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n254), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n261), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n268) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_U46 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n257), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n251) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_U45 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n266), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n252), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n265), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n241), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n254), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n243) );
  AND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_U44 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n266), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n252), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n241) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_U43 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n275), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n257), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n265) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_U42 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n264), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n281), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n252) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_U41 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n261), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n264) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_U40 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n272), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n273), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n266) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_U39 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n273), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n254), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n262) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_U38 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n271), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n273) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_U37 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n275), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n281), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n260) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_U36 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n258), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n275) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_U35 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n258), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n240), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n261), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n240), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n254), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n245) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_U34 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n239), .B(
        Red_StateRegOutput[14]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n254) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_U33 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n238), .B(
        F_SD2_RedSB_inst_n26), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n239) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_U32 ( .A(
        Red_StateRegOutput[16]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n238), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n261) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_U31 ( .A(
        F_SD2_RedSB_inst_n27), .B(F_SD2_RedSB_inst_n25), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n238) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_U30 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n257), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n281), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n271), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n240) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_U29 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n237), .B(
        Red_StateRegOutput[17]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n271) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_U28 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n236), .B(
        F_SD2_RedSB_inst_n26), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n281) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_U27 ( .A(
        Red_StateRegOutput[19]), .B(F_SD2_RedSB_inst_n28), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n236) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_U26 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n235), .B(
        Red_StateRegOutput[15]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n257) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_U25 ( .A(
        F_SD2_RedSB_inst_n26), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n237), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n235) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_U24 ( .A(
        F_SD2_RedSB_inst_n25), .B(F_SD2_RedSB_inst_n28), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n237) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_U23 ( .A(
        Red_StateRegOutput[20]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n234), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n258) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_U22 ( .A(
        F_SD2_RedSB_inst_n27), .B(F_SD2_RedSB_inst_n28), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n234) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_U21 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n233), .B(
        Red_StateRegOutput[18]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n272) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_U20 ( .A(
        F_SD2_RedSB_inst_n27), .B(F_SD2_RedSB_inst_n26), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n233) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_U19 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n217), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n221), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n227), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n231), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n232), .ZN(Red_Feedback[95])
         );
  NOR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_U18 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n221), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n231), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n227), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n232) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_U17 ( .A(
        Red_StateRegOutput[19]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n230), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n231) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_U16 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n285), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n286), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n228), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n229), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n230) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_U15 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n279), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n280), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n278), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n229) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_U14 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n284), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n282), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n284), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n283), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n281), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n228) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_U13 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n225), .B2(
        Red_StateRegOutput[16]), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n226), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n227) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_U12 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n225), .B2(
        Red_StateRegOutput[16]), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n217), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n226) );
  AOI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_U11 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n271), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n222), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n223), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n224), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n225) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_U10 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n262), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n286), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n271), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n263), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n224) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_U9 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n270), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n269), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n267), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n268), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n223) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_U8 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n285), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n259), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n276), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n222) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_U7 ( .A(
        Red_StateRegOutput[15]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n220), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n221) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_U6 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n218), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n219), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n220) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_U5 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n265), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n256), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n282), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n274), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n219) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_U4 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n251), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n250), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n249), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n218) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_U3 ( .A(
        Red_StateRegOutput[14]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n246), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_18_n217) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_U73 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n284), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n283), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n282), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n281), .ZN(Red_Feedback[96])
         );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_U72 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n280), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n281), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n279), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n283) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_U71 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n280), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n281), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n282), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n279) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_U70 ( .A(
        Red_StateRegOutput[19]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n278), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n282) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_U69 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n277), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n276), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n278) );
  NAND4_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_U68 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n275), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n274), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n273), .A4(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n272), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n276) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_U67 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n271), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n270), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n269), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n268), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n277) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_U66 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n267), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n268) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_U65 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n274), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n266), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n265), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n264), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n270) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_U64 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n263), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n265) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_U63 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n262), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n272), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n261), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n260), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n266) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_U62 ( .A(
        Red_StateRegOutput[15]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n259), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n281) );
  NOR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_U61 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n258), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n257), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n256), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n259) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_U60 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n255), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n254), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n255), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n253), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n252), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n256) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_U59 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n273), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n263), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n252) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_U58 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n251), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n250), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n263) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_U57 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n275), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n262), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n253) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_U56 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n271), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n269), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n254) );
  AOI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_U55 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n275), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n249), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n248), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n247), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n257) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_U54 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n246), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n245), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n275), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n247) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_U53 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n271), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n244), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n249) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_U52 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n245), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n271) );
  NOR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_U51 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n251), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n244), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n250), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n258) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_U50 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n260), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n248), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n250) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_U49 ( .A(
        Red_StateRegOutput[14]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n243), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n280) );
  AOI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_U48 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n275), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n242), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n241), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n240), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n243) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_U47 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n251), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n239), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n255), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n238), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n240) );
  OR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_U46 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n251), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n239), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n260), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n238) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_U45 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n237), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n248), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n244), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n255) );
  NOR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_U44 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n237), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n236), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n272), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n241) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_U43 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n274), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n262), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n246), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n235), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n236) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_U42 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n234), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n260), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n233), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n242) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_U41 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n232), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n246), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n262), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n233) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_U40 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n231), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n234) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_U39 ( .A(
        Red_StateRegOutput[16]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n230), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n284) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_U38 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n262), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n229), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n228), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n230) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_U37 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n267), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n227), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n226), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n264), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n228) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_U36 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n244), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n225), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n264) );
  NAND4_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_U35 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n237), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n269), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n274), .A4(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n227), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n226) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_U34 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n272), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n269) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_U33 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n237), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n273), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n262), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n231), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n267) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_U32 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n245), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n248), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n231) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_U31 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n244), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n239), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n273) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_U30 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n245), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n225), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n239) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_U29 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n260), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n237) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_U28 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n274), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n224), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n223), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n251), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n229) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_U27 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n232), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n244), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n261), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n244), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n235), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n224) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_U26 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n275), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n245), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n235) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_U25 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n227), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n275) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_U24 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n251), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n261) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_U23 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n227), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n272), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n251) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_U22 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n222), .B(
        Red_StateRegOutput[18]), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n272) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_U21 ( .A(
        F_SD2_RedSB_inst_n26), .B(F_SD2_RedSB_inst_n27), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n222) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_U20 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n221), .B(
        Red_StateRegOutput[17]), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n227) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_U19 ( .A(
        F_SD2_RedSB_inst_n25), .B(F_SD2_RedSB_inst_n28), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n221) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_U18 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n246), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n244) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_U17 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n220), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n219), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n246) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_U16 ( .A(
        F_SD2_RedSB_inst_n28), .B(Red_StateRegOutput[15]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n220) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_U15 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n223), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n232) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_U14 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n260), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n245), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n223) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_U13 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n218), .B(
        Red_StateRegOutput[19]), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n245) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_U12 ( .A(
        F_SD2_RedSB_inst_n26), .B(F_SD2_RedSB_inst_n28), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n218) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_U11 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n217), .B(
        F_SD2_RedSB_inst_n27), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n260) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_U10 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n219), .B(
        Red_StateRegOutput[14]), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n217) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_U9 ( .A(
        F_SD2_RedSB_inst_n25), .B(F_SD2_RedSB_inst_n26), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n219) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_U8 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n248), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n274) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_U7 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n216), .B(
        Red_StateRegOutput[20]), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n248) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_U6 ( .A(
        F_SD2_RedSB_inst_n27), .B(F_SD2_RedSB_inst_n28), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n216) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_U5 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n225), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n262) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_U4 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n215), .B(
        F_SD2_RedSB_inst_n27), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n225) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_U3 ( .A(
        Red_StateRegOutput[16]), .B(F_SD2_RedSB_inst_n25), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_19_n215) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_U65 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n283), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n282), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n281), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n280), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n279), .ZN(Red_Feedback[97])
         );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_U64 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n283), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n282), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n281), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n279) );
  MUX2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_U63 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n283), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n282), .S(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n278), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n280) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_U62 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n277), .B(
        Red_StateRegOutput[16]), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n278) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_U61 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n276), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n275), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n274), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n277) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_U60 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n273), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n274) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_U59 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n272), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n271), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n270), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n269), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n268), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n273) );
  AND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_U58 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n267), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n266), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n265), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n269) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_U57 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n266), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n264), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n263), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n262), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n275) );
  AOI222_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_U56 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n261), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n260), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n261), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n259), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n260), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n259), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n263) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_U55 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n258), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n268), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n259) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_U54 ( .A(
        Red_StateRegOutput[14]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n257), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n281) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_U53 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n268), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n256), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n255), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n257) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_U52 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n268), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n254), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n262), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n255) );
  AOI222_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_U51 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n261), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n260), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n261), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n253), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n260), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n253), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n254) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_U50 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n276), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n258), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n253) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_U49 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n252), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n251), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n250), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n249), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n256) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_U48 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n276), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n266), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n248), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n247), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n252) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_U47 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n264), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n247) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_U46 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n272), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n258), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n264) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_U45 ( .A(
        Red_StateRegOutput[15]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n246), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n282) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_U44 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n248), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n262), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n245), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n244), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n246) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_U43 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n248), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n243), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n244) );
  AOI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_U42 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n271), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n242), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n241), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n240), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n245) );
  NOR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_U41 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n270), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n239), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n250), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n240) );
  AND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_U40 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n238), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n268), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n260), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n241) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_U39 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n248), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n266), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n260) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_U38 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n251), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n237), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n249), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n238) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_U37 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n276), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n270), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n249) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_U36 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n258), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n236), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n262) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_U35 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n237), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n258) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_U34 ( .A(
        Red_StateRegOutput[19]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n235), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n283) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_U33 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n234), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n237), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n233), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n237), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n232), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n235) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_U32 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n251), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n268), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n267), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n236), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n271), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n232) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_U31 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n250), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n276), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n271) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_U30 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n237), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n248), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n250) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_U29 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n239), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n272), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n236) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_U28 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n242), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n265), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n243), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n233) );
  AND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_U27 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n261), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n231), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n243) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_U26 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n276), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n248), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n265) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_U25 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n230), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n229), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n248) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_U24 ( .A(
        F_SD2_RedSB_inst_n25), .B(Red_StateRegOutput[15]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n230) );
  OR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_U23 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n261), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n231), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n242) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_U22 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n268), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n266), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n231) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_U21 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n228), .B(
        Red_StateRegOutput[14]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n268) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_U20 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n227), .B(
        F_SD2_RedSB_inst_n26), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n228) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_U19 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n267), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n270), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n261) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_U18 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n272), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n270) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_U17 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n226), .B(
        Red_StateRegOutput[17]), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n272) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_U16 ( .A(
        F_SD2_RedSB_inst_n25), .B(F_SD2_RedSB_inst_n28), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n226) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_U15 ( .A(
        Red_StateRegOutput[19]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n229), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n237) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_U14 ( .A(
        F_SD2_RedSB_inst_n28), .B(F_SD2_RedSB_inst_n26), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n229) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_U13 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n225), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n234) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_U12 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n267), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n239), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n224), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n225) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_U11 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n267), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n239), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n276), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n224) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_U10 ( .A(
        Red_StateRegOutput[16]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n227), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n276) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_U9 ( .A(
        F_SD2_RedSB_inst_n27), .B(F_SD2_RedSB_inst_n25), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n227) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_U8 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n266), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n239) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_U7 ( .A(
        Red_StateRegOutput[20]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n223), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n266) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_U6 ( .A(
        F_SD2_RedSB_inst_n27), .B(F_SD2_RedSB_inst_n28), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n223) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_U5 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n251), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n267) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_U4 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n222), .B(
        Red_StateRegOutput[18]), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n251) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_U3 ( .A(
        F_SD2_RedSB_inst_n27), .B(F_SD2_RedSB_inst_n26), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_20_n222) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_U69 ( .A(
        Red_StateRegOutput[22]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n280), .Z(Red_Feedback[98])
         );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_U68 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n279), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n278), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n280) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_U67 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n277), .B2(
        Red_StateRegOutput[23]), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n276), .C2(
        Red_StateRegOutput[26]), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n275), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n278) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_U66 ( .A1(
        Red_StateRegOutput[23]), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n277), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n276), .B2(
        Red_StateRegOutput[26]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n275) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_U65 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n274), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n273), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n276) );
  AOI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_U64 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n272), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n271), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n270), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n269), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n273) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_U63 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n268), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n267), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n266), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n265), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n264), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n269) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_U62 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n268), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n263), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n262), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n270) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_U61 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n268), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n263), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n261), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n262) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_U60 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n260), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n259), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n258), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n271) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_U59 ( .A(
        Red_StateRegOutput[21]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n257), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n274) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_U58 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n244), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n243), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n245), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n242), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n241), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n277) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_U57 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n240), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n239), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n238), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n241) );
  AOI222_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_U56 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n255), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n253), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n255), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n237), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n253), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n237), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n239) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_U55 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n247), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n267), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n237) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_U54 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n263), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n251), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n253) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_U53 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n236), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n255) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_U52 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n256), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n235), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n242) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_U51 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n261), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n263), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n234), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n243) );
  NOR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_U50 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n267), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n249), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n259), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n234) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_U49 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n250), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n251), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n259) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_U48 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n268), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n233), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n249) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_U47 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n256), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n267) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_U46 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n247), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n250), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n261) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_U45 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n264), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n260), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n232), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n279) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_U44 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n251), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n231), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n230), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n232) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_U43 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n251), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n229), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n252), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n230) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_U42 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n240), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n252) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_U41 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n247), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n265), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n240) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_U40 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n244), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n233), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n265) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_U39 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n246), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n248), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n256), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n263), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n229) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_U38 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n245), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n250), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n248) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_U37 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n266), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n247), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n246) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_U36 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n272), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n228), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n258), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n231) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_U35 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n236), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n227), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n258) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_U34 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n245), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n233), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n228) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_U33 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n236), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n227), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n260) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_U32 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n233), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n256), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n227) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_U31 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n226), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n225), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n256) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_U30 ( .A(
        Red_StateRegOutput[21]), .B(F_SD2_RedSB_inst_n29), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n226) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_U29 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n263), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n233) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_U28 ( .A(
        Red_StateRegOutput[27]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n224), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n263) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_U27 ( .A(
        F_SD2_RedSB_inst_n32), .B(F_SD2_RedSB_inst_n31), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n224) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_U26 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n244), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n268), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n236) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_U25 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n266), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n268) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_U24 ( .A(
        Red_StateRegOutput[25]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n225), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n266) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_U23 ( .A(
        F_SD2_RedSB_inst_n30), .B(F_SD2_RedSB_inst_n31), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n225) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_U22 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n245), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n244) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_U21 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n223), .B(
        Red_StateRegOutput[24]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n245) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_U20 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n235), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n264) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_U19 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n254), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n251), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n235) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_U18 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n222), .B(
        F_SD2_RedSB_inst_n30), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n251) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_U17 ( .A(
        Red_StateRegOutput[22]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n223), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n222) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_U16 ( .A(
        F_SD2_RedSB_inst_n32), .B(F_SD2_RedSB_inst_n29), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n223) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_U15 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n247), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n250), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n254) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_U14 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n238), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n250) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_U13 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n221), .B(
        Red_StateRegOutput[23]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n238) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_U12 ( .A(
        F_SD2_RedSB_inst_n29), .B(F_SD2_RedSB_inst_n31), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n221) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_U11 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n272), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n247) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_U10 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n220), .B(
        F_SD2_RedSB_inst_n30), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n272) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_U9 ( .A(
        Red_StateRegOutput[26]), .B(F_SD2_RedSB_inst_n32), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n220) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_U8 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n215), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n217), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n256), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n219), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n257) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_U7 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n251), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n218), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n250), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n249), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n219) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_U6 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n247), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n248), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n245), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n246), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n218) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_U5 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n254), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n255), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n252), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n216), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n217) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_U4 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n267), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n216) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_U3 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n255), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n254), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n253), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_21_n215) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_U68 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n273), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n274) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_U67 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n272), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n271), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n275) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_U66 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n267), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n266), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n269) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_U65 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n272), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n271), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n264), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n265) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_U64 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n260), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n259), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n267), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n268), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n261) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_U63 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n258), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n257), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n268) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_U62 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n256), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n267), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n255), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n254), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n260) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_U61 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n253), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n267) );
  NOR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_U60 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n252), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n251), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n250), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n262) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_U59 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n270), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n263) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_U58 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n258), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n257), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n270) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_U57 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n272), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n249), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n257) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_U56 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n252), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n273), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n246) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_U55 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n264), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n250), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n273) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_U54 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n253), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n259), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n250) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_U53 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n266), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n264) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_U52 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n252), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n259), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n248) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_U51 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n278), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n259) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_U50 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n278), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n249), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n245) );
  AND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_U49 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n277), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n271), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n258) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_U48 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n272), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n253), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n255) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_U47 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n251), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n272) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_U46 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n251), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n277), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n256) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_U45 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n252), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n277) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_U44 ( .A(
        Red_StateRegOutput[26]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n244), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n278) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_U43 ( .A(
        F_SD2_RedSB_inst_n31), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n243), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n266) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_U42 ( .A(
        Red_StateRegOutput[23]), .B(F_SD2_RedSB_inst_n29), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n243) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_U41 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n254), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n276) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_U40 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n271), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n247), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n254) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_U39 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n249), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n247) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_U38 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n242), .B(
        Red_StateRegOutput[21]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n249) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_U37 ( .A(
        F_SD2_RedSB_inst_n29), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n241), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n242) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_U36 ( .A(
        Red_StateRegOutput[25]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n241), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n271) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_U35 ( .A(
        F_SD2_RedSB_inst_n31), .B(F_SD2_RedSB_inst_n30), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n241) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_U34 ( .A(
        Red_StateRegOutput[27]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n240), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n251) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_U33 ( .A(
        F_SD2_RedSB_inst_n31), .B(F_SD2_RedSB_inst_n32), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n240) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_U32 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n239), .B(
        Red_StateRegOutput[24]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n252) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_U31 ( .A(
        F_SD2_RedSB_inst_n29), .B(F_SD2_RedSB_inst_n32), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n239) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_U30 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n238), .B(
        Red_StateRegOutput[22]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n253) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_U29 ( .A(
        F_SD2_RedSB_inst_n29), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n244), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n238) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_U28 ( .A(
        F_SD2_RedSB_inst_n30), .B(F_SD2_RedSB_inst_n32), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n244) );
  AOI222_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_U27 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n221), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n228), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n221), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n233), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n228), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n237), .ZN(Red_Feedback[99])
         );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_U26 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n236), .B(
        Red_StateRegOutput[22]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n237) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_U25 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n234), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n235), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n236) );
  AOI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_U24 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n273), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n263), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n261), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n262), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n235) );
  NAND4_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_U23 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n249), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n252), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n264), .A4(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n255), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n234) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_U22 ( .A(
        Red_StateRegOutput[26]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n232), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n233) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_U21 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n229), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n278), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n230), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n278), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n231), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n232) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_U20 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n277), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n276), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n275), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n276), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n274), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n231) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_U19 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n270), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n269), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n268), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n230) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_U18 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n272), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n271), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n265), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n229) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_U17 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n227), .B(
        Red_StateRegOutput[23]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n228) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_U16 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n266), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n222), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n226), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n227) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_U15 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n247), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n246), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n225), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n226) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_U14 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n224), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n255), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n224), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n245), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n264), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n225) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_U13 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n217), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n223), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n224) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_U12 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n251), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n248), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n258), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n245), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n223) );
  NOR4_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_U11 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n251), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n252), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n253), .A4(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n276), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n222) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_U10 ( .A(
        Red_StateRegOutput[21]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n220), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n221) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_U9 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n249), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n216), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n219), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n220) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_U8 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n249), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n217), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n218), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n219) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_U7 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n258), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n255), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n259), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n266), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n218) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_U6 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n278), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n256), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n258), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n255), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n217) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_U5 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n250), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n214), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n271), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n215), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n216) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_U4 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n264), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n272), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n253), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n248), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n215) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_U3 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n252), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n264), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_22_n214) );
  MUX2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_U54 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n240), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n239), .S(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n238), .Z(Red_Feedback[100])
         );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_U53 ( .A(
        Red_StateRegOutput[23]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n237), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n238) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_U52 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n236), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n235), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n234), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n233), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n237) );
  OR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_U51 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n232), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n231), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n230), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n233) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_U50 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n229), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n228), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n227), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n234) );
  AOI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_U49 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n226), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n225), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n224), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n223), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n236) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_U48 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n222), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n221), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n220), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n221), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n219), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n223) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_U47 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n226), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n225), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n218), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n221) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_U46 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n217), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n216), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n225) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_U45 ( .A(
        Red_StateRegOutput[26]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n215), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n239) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_U44 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n214), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n230), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n213), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n212), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n215) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_U43 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n228), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n226), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n211), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n232), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n212) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_U42 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n210), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n228), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n210), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n226), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n216), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n213) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_U41 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n220), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n216) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_U40 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n209), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n226) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_U39 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n208), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n207), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n228) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_U38 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n219), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n206), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n205), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n210) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_U37 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n219), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n206), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n208), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n205) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_U36 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n235), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n208) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_U35 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n222), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n204), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n229), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n214) );
  AND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_U34 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n206), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n219), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n204) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_U33 ( .A(
        Red_StateRegOutput[22]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n203), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n240) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_U32 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n202), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n201), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n200), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n201), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n199), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n203) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_U31 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n198), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n197), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n230), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n209), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n199) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_U30 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n227), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n220), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n218), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n197) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_U29 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n207), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n218) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_U28 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n222), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n201), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n227) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_U27 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n198), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n230), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n209), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n230), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n217), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n200) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_U26 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n231), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n206), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n209) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_U25 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n207), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n235), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n220), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n230) );
  AOI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_U24 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n229), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n211), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n207), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n224), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n198) );
  NOR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_U23 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n231), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n220), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n201), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n224) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_U22 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n219), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n220), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n211) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_U21 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n196), .B(
        Red_StateRegOutput[26]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n220) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_U20 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n201), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n219) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_U19 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n232), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n206), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n229) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_U18 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n195), .B(
        Red_StateRegOutput[25]), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n206) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_U17 ( .A(
        F_SD2_RedSB_inst_n31), .B(F_SD2_RedSB_inst_n30), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n195) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_U16 ( .A(
        Red_StateRegOutput[27]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n194), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n201) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_U15 ( .A(
        F_SD2_RedSB_inst_n31), .B(F_SD2_RedSB_inst_n32), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n194) );
  NOR4_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_U14 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n207), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n231), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n232), .A4(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n235), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n202) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_U13 ( .A(
        Red_StateRegOutput[23]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n193), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n235) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_U12 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n217), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n232) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_U11 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n192), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n193), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n217) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_U10 ( .A(
        F_SD2_RedSB_inst_n29), .B(F_SD2_RedSB_inst_n31), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n193) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_U9 ( .A(
        F_SD2_RedSB_inst_n30), .B(Red_StateRegOutput[21]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n192) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_U8 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n222), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n231) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_U7 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n191), .B(
        Red_StateRegOutput[24]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n222) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_U6 ( .A(
        F_SD2_RedSB_inst_n29), .B(F_SD2_RedSB_inst_n32), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n191) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_U5 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n190), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n196), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n207) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_U4 ( .A(
        F_SD2_RedSB_inst_n30), .B(F_SD2_RedSB_inst_n32), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n196) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_U3 ( .A(
        F_SD2_RedSB_inst_n29), .B(Red_StateRegOutput[22]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_23_n190) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_U70 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n290), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n289), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n288), .ZN(Red_Feedback[101])
         );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_U69 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n290), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n287), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n288) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_U68 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n286), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n285), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n284), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n287) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_U67 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n283), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n282), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n286), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n284) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_U66 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n289), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n285) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_U65 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n283), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n282), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n281), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n289) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_U64 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n282), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n286), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n283), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n281) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_U63 ( .A(
        Red_StateRegOutput[26]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n268), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n282) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_U62 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n267), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n266), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n265), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n269), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n268) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_U61 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n264), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n274), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n263), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n262), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n261), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n265) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_U60 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n260), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n259), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n278), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n258), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n263) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_U59 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n262), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n274) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_U58 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n273), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n272), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n264) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_U57 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n257), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n266) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_U56 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n256), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n255), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n254), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n267) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_U55 ( .A(
        Red_StateRegOutput[23]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n253), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n283) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_U54 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n252), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n262), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n251), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n250), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n253) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_U53 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n278), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n257), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n249), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n250) );
  NAND4_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_U52 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n254), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n248), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n276), .A4(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n262), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n251) );
  AOI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_U51 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n271), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n247), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n246), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n277), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n252) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_U50 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n258), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n259), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n245), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n277) );
  NOR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_U49 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n278), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n244), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n280), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n246) );
  AND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_U48 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n258), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n259), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n280) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_U47 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n243), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n259) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_U46 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n249), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n269), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n271) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_U45 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n276), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n279), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n257) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_U44 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n262), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n269), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n279) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_U43 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n244), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n256), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n245) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_U42 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n241), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n247), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n256) );
  AND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_U41 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n243), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n242), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n261) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_U40 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n278), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n272), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n242) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_U39 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n249), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n273), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n243) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_U38 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n255), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n273) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_U37 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n249), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n247), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n248) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_U36 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n275), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n255), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n254) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_U35 ( .A(
        Red_StateRegOutput[25]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n240), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n255) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_U34 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n278), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n275) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_U33 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n269), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n244) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_U32 ( .A(
        Red_StateRegOutput[26]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n239), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n269) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_U31 ( .A(
        F_SD2_RedSB_inst_n30), .B(F_SD2_RedSB_inst_n32), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n239) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_U30 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n262), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n241), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n270) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_U29 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n249), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n241) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_U28 ( .A(
        Red_StateRegOutput[24]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n238), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n249) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_U27 ( .A(
        F_SD2_RedSB_inst_n29), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n237), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n262) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_U26 ( .A(
        Red_StateRegOutput[23]), .B(F_SD2_RedSB_inst_n31), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n237) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_U25 ( .A(
        F_SD2_RedSB_inst_n30), .B(F_SD2_RedSB_inst_n31), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n240) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_U24 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n276), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n247), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n258) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_U23 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n272), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n247) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_U22 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n236), .B(
        Red_StateRegOutput[27]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n272) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_U21 ( .A(
        F_SD2_RedSB_inst_n31), .B(F_SD2_RedSB_inst_n32), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n236) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_U20 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n260), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n276) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_U19 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n235), .B(
        Red_StateRegOutput[22]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n260) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_U18 ( .A(
        F_SD2_RedSB_inst_n30), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n238), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n235) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_U17 ( .A(
        F_SD2_RedSB_inst_n29), .B(F_SD2_RedSB_inst_n32), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n238) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_U16 ( .A(
        Red_StateRegOutput[22]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n234), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n290) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_U15 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n258), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n230), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n232), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n233), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n234) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_U14 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n261), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n269), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n261), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n248), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n260), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n233) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_U13 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n243), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n257), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n242), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n257), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n231), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n232) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_U12 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n260), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n245), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n231) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_U11 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n278), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n270), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n244), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n254), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n230) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_U10 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n229), .B(
        Red_StateRegOutput[21]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n286) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_U9 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n225), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n277), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n228), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n229) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_U8 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n276), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n226), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n275), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n227), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n228) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_U7 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n274), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n272), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n273), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n227) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_U6 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n269), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n270), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n273), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n271), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n226) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_U5 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n280), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n279), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n278), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n225) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_U4 ( .A(
        Red_StateRegOutput[21]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n224), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n278) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_U3 ( .A(
        F_SD2_RedSB_inst_n29), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n240), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_24_n224) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_U73 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n277), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n276), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n279), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n278) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_U72 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n275), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n274), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n273), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n277) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_U71 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n272), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n279) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_U70 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n266), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n265), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n264), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n267) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_U69 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n265), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n269) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_U68 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n280), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n263) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_U67 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n261), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n260), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n280) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_U66 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n264), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n281), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n258), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n276) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_U65 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n283), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n275), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n259) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_U64 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n264), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n257), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n283) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_U63 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n261), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n262), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n255), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n285), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n256) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_U62 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n272), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n254), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n285) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_U61 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n270), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n253), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n282) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_U60 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n286), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n274) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_U59 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n257), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n252), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n286) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_U58 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n260), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n271), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n251), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n249) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_U57 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n273), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n248), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n247), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n250) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_U56 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n284), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n247) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_U55 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n270), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n253), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n284) );
  OR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_U54 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n275), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n254), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n253) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_U53 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n266), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n270) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_U52 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n255), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n275), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n248) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_U51 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n281), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n255) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_U50 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n272), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n245), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n244), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n246) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_U49 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n260), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n262), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n243), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n242), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n244) );
  OR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_U48 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n251), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n271), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n268), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n242) );
  OR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_U47 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n281), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n254), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n261), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n268) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_U46 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n257), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n251) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_U45 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n266), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n252), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n265), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n241), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n254), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n243) );
  AND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_U44 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n266), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n252), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n241) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_U43 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n275), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n257), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n265) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_U42 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n264), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n281), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n252) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_U41 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n261), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n264) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_U40 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n272), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n273), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n266) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_U39 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n273), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n254), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n262) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_U38 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n271), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n273) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_U37 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n275), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n281), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n260) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_U36 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n258), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n275) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_U35 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n258), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n240), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n261), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n240), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n254), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n245) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_U34 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n239), .B(
        Red_StateRegOutput[21]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n254) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_U33 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n238), .B(
        F_SD2_RedSB_inst_n30), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n239) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_U32 ( .A(
        Red_StateRegOutput[23]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n238), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n261) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_U31 ( .A(
        F_SD2_RedSB_inst_n31), .B(F_SD2_RedSB_inst_n29), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n238) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_U30 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n257), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n281), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n271), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n240) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_U29 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n237), .B(
        Red_StateRegOutput[24]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n271) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_U28 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n236), .B(
        F_SD2_RedSB_inst_n30), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n281) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_U27 ( .A(
        Red_StateRegOutput[26]), .B(F_SD2_RedSB_inst_n32), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n236) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_U26 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n235), .B(
        Red_StateRegOutput[22]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n257) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_U25 ( .A(
        F_SD2_RedSB_inst_n30), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n237), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n235) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_U24 ( .A(
        F_SD2_RedSB_inst_n29), .B(F_SD2_RedSB_inst_n32), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n237) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_U23 ( .A(
        Red_StateRegOutput[27]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n234), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n258) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_U22 ( .A(
        F_SD2_RedSB_inst_n31), .B(F_SD2_RedSB_inst_n32), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n234) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_U21 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n233), .B(
        Red_StateRegOutput[25]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n272) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_U20 ( .A(
        F_SD2_RedSB_inst_n31), .B(F_SD2_RedSB_inst_n30), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n233) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_U19 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n217), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n221), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n227), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n231), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n232), .ZN(Red_Feedback[102])
         );
  NOR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_U18 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n221), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n231), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n227), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n232) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_U17 ( .A(
        Red_StateRegOutput[26]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n230), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n231) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_U16 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n285), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n286), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n228), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n229), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n230) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_U15 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n279), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n280), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n278), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n229) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_U14 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n284), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n282), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n284), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n283), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n281), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n228) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_U13 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n225), .B2(
        Red_StateRegOutput[23]), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n226), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n227) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_U12 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n225), .B2(
        Red_StateRegOutput[23]), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n217), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n226) );
  AOI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_U11 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n271), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n222), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n223), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n224), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n225) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_U10 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n262), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n286), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n271), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n263), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n224) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_U9 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n270), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n269), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n267), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n268), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n223) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_U8 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n285), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n259), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n276), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n222) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_U7 ( .A(
        Red_StateRegOutput[22]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n220), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n221) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_U6 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n218), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n219), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n220) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_U5 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n265), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n256), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n282), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n274), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n219) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_U4 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n251), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n250), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n249), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n218) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_U3 ( .A(
        Red_StateRegOutput[21]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n246), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_25_n217) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_U73 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n284), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n283), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n282), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n281), .ZN(Red_Feedback[103])
         );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_U72 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n280), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n281), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n279), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n283) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_U71 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n280), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n281), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n282), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n279) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_U70 ( .A(
        Red_StateRegOutput[26]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n278), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n282) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_U69 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n277), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n276), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n278) );
  NAND4_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_U68 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n275), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n274), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n273), .A4(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n272), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n276) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_U67 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n271), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n270), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n269), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n268), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n277) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_U66 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n267), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n268) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_U65 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n274), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n266), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n265), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n264), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n270) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_U64 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n263), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n265) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_U63 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n262), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n272), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n261), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n260), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n266) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_U62 ( .A(
        Red_StateRegOutput[22]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n259), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n281) );
  NOR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_U61 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n258), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n257), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n256), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n259) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_U60 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n255), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n254), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n255), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n253), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n252), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n256) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_U59 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n273), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n263), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n252) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_U58 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n251), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n250), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n263) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_U57 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n275), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n262), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n253) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_U56 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n271), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n269), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n254) );
  AOI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_U55 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n275), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n249), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n248), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n247), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n257) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_U54 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n246), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n245), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n275), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n247) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_U53 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n271), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n244), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n249) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_U52 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n245), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n271) );
  NOR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_U51 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n251), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n244), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n250), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n258) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_U50 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n260), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n248), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n250) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_U49 ( .A(
        Red_StateRegOutput[21]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n243), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n280) );
  AOI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_U48 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n275), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n242), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n241), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n240), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n243) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_U47 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n251), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n239), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n255), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n238), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n240) );
  OR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_U46 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n251), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n239), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n260), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n238) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_U45 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n237), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n248), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n244), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n255) );
  NOR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_U44 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n237), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n236), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n272), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n241) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_U43 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n274), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n262), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n246), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n235), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n236) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_U42 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n234), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n260), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n233), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n242) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_U41 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n232), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n246), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n262), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n233) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_U40 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n231), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n234) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_U39 ( .A(
        Red_StateRegOutput[23]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n230), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n284) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_U38 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n262), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n229), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n228), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n230) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_U37 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n267), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n227), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n226), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n264), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n228) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_U36 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n244), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n225), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n264) );
  NAND4_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_U35 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n237), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n269), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n274), .A4(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n227), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n226) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_U34 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n272), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n269) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_U33 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n237), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n273), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n262), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n231), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n267) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_U32 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n245), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n248), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n231) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_U31 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n244), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n239), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n273) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_U30 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n245), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n225), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n239) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_U29 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n260), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n237) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_U28 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n274), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n224), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n223), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n251), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n229) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_U27 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n232), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n244), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n261), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n244), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n235), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n224) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_U26 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n275), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n245), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n235) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_U25 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n227), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n275) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_U24 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n251), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n261) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_U23 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n227), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n272), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n251) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_U22 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n222), .B(
        Red_StateRegOutput[25]), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n272) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_U21 ( .A(
        F_SD2_RedSB_inst_n30), .B(F_SD2_RedSB_inst_n31), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n222) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_U20 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n221), .B(
        Red_StateRegOutput[24]), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n227) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_U19 ( .A(
        F_SD2_RedSB_inst_n29), .B(F_SD2_RedSB_inst_n32), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n221) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_U18 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n246), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n244) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_U17 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n220), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n219), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n246) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_U16 ( .A(
        F_SD2_RedSB_inst_n32), .B(Red_StateRegOutput[22]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n220) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_U15 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n223), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n232) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_U14 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n260), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n245), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n223) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_U13 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n218), .B(
        Red_StateRegOutput[26]), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n245) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_U12 ( .A(
        F_SD2_RedSB_inst_n30), .B(F_SD2_RedSB_inst_n32), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n218) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_U11 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n217), .B(
        F_SD2_RedSB_inst_n31), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n260) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_U10 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n219), .B(
        Red_StateRegOutput[21]), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n217) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_U9 ( .A(
        F_SD2_RedSB_inst_n29), .B(F_SD2_RedSB_inst_n30), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n219) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_U8 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n248), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n274) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_U7 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n216), .B(
        Red_StateRegOutput[27]), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n248) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_U6 ( .A(
        F_SD2_RedSB_inst_n31), .B(F_SD2_RedSB_inst_n32), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n216) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_U5 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n225), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n262) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_U4 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n215), .B(
        F_SD2_RedSB_inst_n31), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n225) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_U3 ( .A(
        Red_StateRegOutput[23]), .B(F_SD2_RedSB_inst_n29), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_26_n215) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_U65 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n283), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n282), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n281), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n280), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n279), .ZN(Red_Feedback[104])
         );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_U64 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n283), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n282), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n281), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n279) );
  MUX2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_U63 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n283), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n282), .S(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n278), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n280) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_U62 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n277), .B(
        Red_StateRegOutput[23]), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n278) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_U61 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n276), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n275), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n274), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n277) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_U60 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n273), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n274) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_U59 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n272), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n271), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n270), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n269), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n268), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n273) );
  AND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_U58 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n267), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n266), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n265), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n269) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_U57 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n266), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n264), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n263), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n262), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n275) );
  AOI222_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_U56 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n261), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n260), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n261), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n259), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n260), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n259), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n263) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_U55 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n258), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n268), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n259) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_U54 ( .A(
        Red_StateRegOutput[21]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n257), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n281) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_U53 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n268), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n256), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n255), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n257) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_U52 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n268), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n254), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n262), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n255) );
  AOI222_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_U51 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n261), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n260), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n261), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n253), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n260), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n253), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n254) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_U50 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n276), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n258), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n253) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_U49 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n252), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n251), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n250), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n249), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n256) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_U48 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n276), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n266), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n248), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n247), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n252) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_U47 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n264), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n247) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_U46 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n272), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n258), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n264) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_U45 ( .A(
        Red_StateRegOutput[22]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n246), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n282) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_U44 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n248), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n262), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n245), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n244), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n246) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_U43 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n248), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n243), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n244) );
  AOI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_U42 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n271), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n242), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n241), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n240), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n245) );
  NOR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_U41 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n270), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n239), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n250), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n240) );
  AND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_U40 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n238), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n268), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n260), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n241) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_U39 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n248), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n266), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n260) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_U38 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n251), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n237), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n249), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n238) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_U37 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n276), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n270), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n249) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_U36 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n258), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n236), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n262) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_U35 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n237), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n258) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_U34 ( .A(
        Red_StateRegOutput[26]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n235), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n283) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_U33 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n234), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n237), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n233), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n237), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n232), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n235) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_U32 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n251), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n268), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n267), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n236), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n271), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n232) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_U31 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n250), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n276), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n271) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_U30 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n237), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n248), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n250) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_U29 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n239), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n272), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n236) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_U28 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n242), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n265), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n243), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n233) );
  AND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_U27 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n261), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n231), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n243) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_U26 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n276), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n248), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n265) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_U25 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n230), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n229), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n248) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_U24 ( .A(
        F_SD2_RedSB_inst_n29), .B(Red_StateRegOutput[22]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n230) );
  OR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_U23 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n261), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n231), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n242) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_U22 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n268), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n266), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n231) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_U21 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n228), .B(
        Red_StateRegOutput[21]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n268) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_U20 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n227), .B(
        F_SD2_RedSB_inst_n30), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n228) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_U19 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n267), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n270), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n261) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_U18 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n272), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n270) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_U17 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n226), .B(
        Red_StateRegOutput[24]), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n272) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_U16 ( .A(
        F_SD2_RedSB_inst_n29), .B(F_SD2_RedSB_inst_n32), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n226) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_U15 ( .A(
        Red_StateRegOutput[26]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n229), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n237) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_U14 ( .A(
        F_SD2_RedSB_inst_n32), .B(F_SD2_RedSB_inst_n30), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n229) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_U13 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n225), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n234) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_U12 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n267), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n239), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n224), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n225) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_U11 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n267), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n239), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n276), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n224) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_U10 ( .A(
        Red_StateRegOutput[23]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n227), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n276) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_U9 ( .A(
        F_SD2_RedSB_inst_n31), .B(F_SD2_RedSB_inst_n29), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n227) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_U8 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n266), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n239) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_U7 ( .A(
        Red_StateRegOutput[27]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n223), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n266) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_U6 ( .A(
        F_SD2_RedSB_inst_n31), .B(F_SD2_RedSB_inst_n32), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n223) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_U5 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n251), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n267) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_U4 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n222), .B(
        Red_StateRegOutput[25]), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n251) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_U3 ( .A(
        F_SD2_RedSB_inst_n31), .B(F_SD2_RedSB_inst_n30), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_27_n222) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_U69 ( .A(
        Red_StateRegOutput[29]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n280), .Z(Red_Feedback[56])
         );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_U68 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n279), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n278), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n280) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_U67 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n277), .B2(
        Red_StateRegOutput[30]), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n276), .C2(
        Red_StateRegOutput[33]), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n275), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n278) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_U66 ( .A1(
        Red_StateRegOutput[30]), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n277), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n276), .B2(
        Red_StateRegOutput[33]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n275) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_U65 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n274), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n273), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n276) );
  AOI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_U64 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n272), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n271), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n270), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n269), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n273) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_U63 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n268), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n267), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n266), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n265), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n264), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n269) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_U62 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n268), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n263), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n262), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n270) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_U61 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n268), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n263), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n261), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n262) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_U60 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n260), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n259), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n258), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n271) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_U59 ( .A(
        Red_StateRegOutput[28]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n257), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n274) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_U58 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n256), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n255), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n254), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n257) );
  OR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_U57 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n267), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n253), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n252), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n254) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_U56 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n251), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n250), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n249), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n252) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_U55 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n250), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n251), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n248), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n253) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_U54 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n247), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n246), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n245), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n244), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n255) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_U53 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n243), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n242), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n241), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n240), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n247) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_U52 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n239), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n238), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n240), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n237), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n236), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n277) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_U51 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n235), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n234), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n233), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n236) );
  AOI222_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_U50 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n251), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n249), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n251), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n232), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n249), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n232), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n234) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_U49 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n242), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n267), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n232) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_U48 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n263), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n246), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n249) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_U47 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n231), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n251) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_U46 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n256), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n230), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n237) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_U45 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n261), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n263), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n229), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n238) );
  NOR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_U44 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n267), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n244), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n259), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n229) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_U43 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n245), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n246), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n259) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_U42 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n268), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n228), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n244) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_U41 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n256), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n267) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_U40 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n242), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n245), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n261) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_U39 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n264), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n260), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n227), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n279) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_U38 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n246), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n226), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n225), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n227) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_U37 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n246), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n224), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n248), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n225) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_U36 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n235), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n248) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_U35 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n242), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n265), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n235) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_U34 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n239), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n228), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n265) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_U33 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n241), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n243), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n256), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n263), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n224) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_U32 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n240), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n245), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n243) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_U31 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n266), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n242), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n241) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_U30 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n272), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n223), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n258), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n226) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_U29 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n231), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n222), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n258) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_U28 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n240), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n228), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n223) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_U27 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n231), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n222), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n260) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_U26 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n228), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n256), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n222) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_U25 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n221), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n220), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n256) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_U24 ( .A(
        Red_StateRegOutput[28]), .B(F_SD2_RedSB_inst_n33), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n221) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_U23 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n263), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n228) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_U22 ( .A(
        Red_StateRegOutput[34]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n219), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n263) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_U21 ( .A(
        F_SD2_RedSB_inst_n36), .B(F_SD2_RedSB_inst_n35), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n219) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_U20 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n239), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n268), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n231) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_U19 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n266), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n268) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_U18 ( .A(
        Red_StateRegOutput[32]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n220), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n266) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_U17 ( .A(
        F_SD2_RedSB_inst_n34), .B(F_SD2_RedSB_inst_n35), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n220) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_U16 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n240), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n239) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_U15 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n218), .B(
        Red_StateRegOutput[31]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n240) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_U14 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n230), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n264) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_U13 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n250), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n246), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n230) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_U12 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n217), .B(
        F_SD2_RedSB_inst_n34), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n246) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_U11 ( .A(
        Red_StateRegOutput[29]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n218), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n217) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_U10 ( .A(
        F_SD2_RedSB_inst_n36), .B(F_SD2_RedSB_inst_n33), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n218) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_U9 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n242), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n245), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n250) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_U8 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n233), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n245) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_U7 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n216), .B(
        Red_StateRegOutput[30]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n233) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_U6 ( .A(
        F_SD2_RedSB_inst_n33), .B(F_SD2_RedSB_inst_n35), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n216) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_U5 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n272), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n242) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_U4 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n215), .B(
        F_SD2_RedSB_inst_n34), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n272) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_U3 ( .A(
        Red_StateRegOutput[33]), .B(F_SD2_RedSB_inst_n36), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_28_n215) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_U67 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n265), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n264), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n270), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n271), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n266) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_U66 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n263), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n262), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n271) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_U65 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n261), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n270), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n260), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n259), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n265) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_U64 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n258), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n270) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_U63 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n272), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n267) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_U62 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n263), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n262), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n272) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_U61 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n274), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n254), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n262) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_U60 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n268), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n255), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n275) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_U59 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n258), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n264), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n255) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_U58 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n269), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n268) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_U57 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n257), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n264), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n253) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_U56 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n277), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n264) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_U55 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n277), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n254), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n251) );
  AND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_U54 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n276), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n273), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n263) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_U53 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n274), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n258), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n260) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_U52 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n256), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n274) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_U51 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n256), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n276), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n261) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_U50 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n257), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n276) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_U49 ( .A(
        Red_StateRegOutput[33]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n250), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n277) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_U48 ( .A(
        F_SD2_RedSB_inst_n35), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n249), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n269) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_U47 ( .A(
        Red_StateRegOutput[30]), .B(F_SD2_RedSB_inst_n33), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n249) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_U46 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n273), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n252), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n259) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_U45 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n254), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n252) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_U44 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n248), .B(
        Red_StateRegOutput[28]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n254) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_U43 ( .A(
        F_SD2_RedSB_inst_n33), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n247), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n248) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_U42 ( .A(
        Red_StateRegOutput[32]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n247), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n273) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_U41 ( .A(
        F_SD2_RedSB_inst_n35), .B(F_SD2_RedSB_inst_n34), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n247) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_U40 ( .A(
        Red_StateRegOutput[34]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n246), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n256) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_U39 ( .A(
        F_SD2_RedSB_inst_n35), .B(F_SD2_RedSB_inst_n36), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n246) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_U38 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n245), .B(
        Red_StateRegOutput[31]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n257) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_U37 ( .A(
        F_SD2_RedSB_inst_n33), .B(F_SD2_RedSB_inst_n36), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n245) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_U36 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n244), .B(
        Red_StateRegOutput[29]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n258) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_U35 ( .A(
        F_SD2_RedSB_inst_n33), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n250), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n244) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_U34 ( .A(
        F_SD2_RedSB_inst_n34), .B(F_SD2_RedSB_inst_n36), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n250) );
  AOI222_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_U33 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n221), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n230), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n221), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n238), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n230), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n243), .ZN(Red_Feedback[57])
         );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_U32 ( .A(
        Red_StateRegOutput[29]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n242), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n243) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_U31 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n255), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n239), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n240), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n241), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n242) );
  NAND4_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_U30 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n254), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n257), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n268), .A4(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n260), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n241) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_U29 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n275), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n267), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n266), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n240) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_U28 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n226), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n239) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_U27 ( .A(
        Red_StateRegOutput[33]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n237), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n238) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_U26 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n277), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n234), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n275), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n236), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n237) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_U25 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n276), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n232), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n235), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n236) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_U24 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n259), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n235) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_U23 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n272), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n231), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n271), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n233), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n234) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_U22 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n273), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n274), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n268), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n232), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n233) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_U21 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n273), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n274), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n232) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_U20 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n270), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n269), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n231) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_U19 ( .A(
        Red_StateRegOutput[30]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n229), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n230) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_U18 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n252), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n222), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n225), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n228), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n229) );
  NAND4_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_U17 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n269), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n259), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n226), .A4(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n227), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n228) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_U16 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n258), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n227) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_U15 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n256), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n257), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n226) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_U14 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n224), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n260), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n224), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n251), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n268), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n225) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_U13 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n217), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n223), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n224) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_U12 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n256), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n253), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n263), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n251), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n223) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_U11 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n257), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n275), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n222) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_U10 ( .A(
        Red_StateRegOutput[28]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n220), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n221) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_U9 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n254), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n216), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n219), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n220) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_U8 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n254), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n217), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n218), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n219) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_U7 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n263), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n260), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n264), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n269), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n218) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_U6 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n277), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n261), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n263), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n260), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n217) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_U5 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n255), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n214), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n273), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n215), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n216) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_U4 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n258), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n253), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n268), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n274), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n215) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_U3 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n257), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n268), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_29_n214) );
  MUX2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_U54 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n240), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n239), .S(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n238), .Z(Red_Feedback[58])
         );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_U53 ( .A(
        Red_StateRegOutput[30]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n237), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n238) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_U52 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n236), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n235), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n234), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n233), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n237) );
  OR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_U51 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n232), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n231), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n230), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n233) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_U50 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n229), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n228), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n227), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n234) );
  AOI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_U49 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n226), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n225), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n224), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n223), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n236) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_U48 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n222), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n221), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n220), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n221), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n219), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n223) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_U47 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n226), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n225), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n218), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n221) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_U46 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n217), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n216), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n225) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_U45 ( .A(
        Red_StateRegOutput[33]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n215), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n239) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_U44 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n214), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n230), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n213), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n212), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n215) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_U43 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n228), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n226), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n211), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n232), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n212) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_U42 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n210), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n228), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n210), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n226), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n216), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n213) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_U41 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n220), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n216) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_U40 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n209), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n226) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_U39 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n208), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n207), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n228) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_U38 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n219), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n206), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n205), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n210) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_U37 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n219), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n206), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n208), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n205) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_U36 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n235), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n208) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_U35 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n222), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n204), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n229), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n214) );
  AND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_U34 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n206), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n219), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n204) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_U33 ( .A(
        Red_StateRegOutput[29]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n203), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n240) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_U32 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n202), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n201), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n200), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n201), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n199), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n203) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_U31 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n198), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n197), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n230), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n209), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n199) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_U30 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n227), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n220), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n218), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n197) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_U29 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n207), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n218) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_U28 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n222), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n201), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n227) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_U27 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n198), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n230), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n209), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n230), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n217), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n200) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_U26 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n231), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n206), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n209) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_U25 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n207), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n235), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n220), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n230) );
  AOI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_U24 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n229), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n211), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n207), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n224), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n198) );
  NOR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_U23 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n231), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n220), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n201), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n224) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_U22 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n219), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n220), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n211) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_U21 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n196), .B(
        Red_StateRegOutput[33]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n220) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_U20 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n201), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n219) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_U19 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n232), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n206), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n229) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_U18 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n195), .B(
        Red_StateRegOutput[32]), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n206) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_U17 ( .A(
        F_SD2_RedSB_inst_n35), .B(F_SD2_RedSB_inst_n34), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n195) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_U16 ( .A(
        Red_StateRegOutput[34]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n194), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n201) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_U15 ( .A(
        F_SD2_RedSB_inst_n35), .B(F_SD2_RedSB_inst_n36), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n194) );
  NOR4_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_U14 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n207), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n231), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n232), .A4(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n235), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n202) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_U13 ( .A(
        Red_StateRegOutput[30]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n193), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n235) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_U12 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n217), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n232) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_U11 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n192), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n193), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n217) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_U10 ( .A(
        F_SD2_RedSB_inst_n33), .B(F_SD2_RedSB_inst_n35), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n193) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_U9 ( .A(
        F_SD2_RedSB_inst_n34), .B(Red_StateRegOutput[28]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n192) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_U8 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n222), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n231) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_U7 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n191), .B(
        Red_StateRegOutput[31]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n222) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_U6 ( .A(
        F_SD2_RedSB_inst_n33), .B(F_SD2_RedSB_inst_n36), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n191) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_U5 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n190), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n196), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n207) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_U4 ( .A(
        F_SD2_RedSB_inst_n34), .B(F_SD2_RedSB_inst_n36), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n196) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_U3 ( .A(
        F_SD2_RedSB_inst_n33), .B(Red_StateRegOutput[29]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_30_n190) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_U71 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n288), .B(
        Red_StateRegOutput[28]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n291) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_U70 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n287), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n286), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n288) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_U69 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n285), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n284), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n283), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n282), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n286) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_U68 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n281), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n282) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_U67 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n280), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n279), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n278), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n277), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n287) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_U66 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n276), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n275), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n274), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n277) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_U65 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n273), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n275), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n272), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n271), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n280) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_U64 ( .A(
        Red_StateRegOutput[33]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n270), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n289) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_U63 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n269), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n268), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n267), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n271), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n270) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_U62 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n266), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n276), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n265), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n264), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n263), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n267) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_U61 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n262), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n261), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n283), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n260), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n265) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_U60 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n264), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n276) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_U59 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n275), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n274), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n266) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_U58 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n259), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n268) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_U57 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n258), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n257), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n256), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n269) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_U56 ( .A(
        Red_StateRegOutput[30]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n255), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n290) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_U55 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n254), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n264), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n253), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n252), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n255) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_U54 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n283), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n259), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n251), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n252) );
  NAND4_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_U53 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n256), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n250), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n279), .A4(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n264), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n253) );
  AOI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_U52 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n273), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n249), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n248), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n281), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n254) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_U51 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n260), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n261), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n247), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n281) );
  NOR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_U50 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n283), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n246), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n285), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n248) );
  AND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_U49 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n260), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n261), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n285) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_U48 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n245), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n261) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_U47 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n251), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n271), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n273) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_U46 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n245), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n243), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n259), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n244) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_U45 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n279), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n284), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n259) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_U44 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n264), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n271), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n284) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_U43 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n246), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n258), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n247) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_U42 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n242), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n249), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n258) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_U41 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n271), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n250), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n263), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n241) );
  AND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_U40 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n245), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n243), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n263) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_U39 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n283), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n274), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n243) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_U38 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n251), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n275), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n245) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_U37 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n257), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n275) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_U36 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n251), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n249), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n250) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_U35 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n278), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n257), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n256) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_U34 ( .A(
        Red_StateRegOutput[32]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n240), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n257) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_U33 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n283), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n278) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_U32 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n271), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n246) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_U31 ( .A(
        Red_StateRegOutput[33]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n239), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n271) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_U30 ( .A(
        F_SD2_RedSB_inst_n34), .B(F_SD2_RedSB_inst_n36), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n239) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_U29 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n264), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n242), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n272) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_U28 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n251), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n242) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_U27 ( .A(
        Red_StateRegOutput[31]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n238), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n251) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_U26 ( .A(
        F_SD2_RedSB_inst_n33), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n237), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n264) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_U25 ( .A(
        Red_StateRegOutput[30]), .B(F_SD2_RedSB_inst_n35), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n237) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_U24 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n236), .B(
        F_SD2_RedSB_inst_n33), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n283) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_U23 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n235), .B(
        Red_StateRegOutput[28]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n236) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_U22 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n240), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n235) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_U21 ( .A(
        F_SD2_RedSB_inst_n34), .B(F_SD2_RedSB_inst_n35), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n240) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_U20 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n279), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n249), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n260) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_U19 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n274), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n249) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_U18 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n234), .B(
        Red_StateRegOutput[34]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n274) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_U17 ( .A(
        F_SD2_RedSB_inst_n35), .B(F_SD2_RedSB_inst_n36), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n234) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_U16 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n262), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n279) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_U15 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n233), .B(
        Red_StateRegOutput[29]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n262) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_U14 ( .A(
        F_SD2_RedSB_inst_n34), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n238), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n233) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_U13 ( .A(
        F_SD2_RedSB_inst_n33), .B(F_SD2_RedSB_inst_n36), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n238) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_U12 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n225), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n229), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n230), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n232), .ZN(Red_Feedback[59])
         );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_U11 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n225), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n231), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n229), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n232) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_U10 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n291), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n231) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_U9 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n290), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n289), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n291), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n230) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_U8 ( .A(
        Red_StateRegOutput[29]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n228), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n229) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_U7 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n260), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n226), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n244), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n227), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n228) );
  MUX2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_U6 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n247), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n241), .S(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n262), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n227) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_U5 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n246), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n256), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n272), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n283), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n226) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_U4 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n290), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n289), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n224), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n225) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_U3 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n289), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n291), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n290), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_31_n224) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_U74 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n287), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n286), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n285), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n284), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n283), .ZN(Red_Feedback[60])
         );
  NOR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_U73 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n286), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n284), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n285), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n283) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_U72 ( .A(
        Red_StateRegOutput[33]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n282), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n284) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_U71 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n281), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n280), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n279), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n278), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n282) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_U70 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n277), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n276), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n277), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n275), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n274), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n278) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_U69 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n273), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n272), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n271), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n279) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_U68 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n270), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n269), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n272), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n271) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_U67 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n268), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n267), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n266), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n270) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_U66 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n265), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n272) );
  AOI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_U65 ( .C1(
        Red_StateRegOutput[30]), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n264), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n263), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n262), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n285) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_U64 ( .A1(
        Red_StateRegOutput[30]), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n264), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n262) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_U63 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n287), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n263) );
  AOI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_U62 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n261), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n260), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n259), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n258), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n264) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_U61 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n257), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n256), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n255), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n254), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n258) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_U60 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n253), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n252), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n251), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n254) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_U59 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n252), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n256) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_U58 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n250), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n261), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n281), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n249), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n259) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_U57 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n273), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n250) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_U56 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n248), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n247), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n273) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_U55 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n280), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n246), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n269), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n260) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_U54 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n251), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n274), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n245), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n269) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_U53 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n276), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n268), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n246) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_U52 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n251), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n244), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n276) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_U51 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n243), .B(
        Red_StateRegOutput[29]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n286) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_U50 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n242), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n241), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n243) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_U49 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n267), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n275), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n252), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n240), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n241) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_U48 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n248), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n249), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n239), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n280), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n240) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_U47 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n265), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n238), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n280) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_U46 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n257), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n237), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n275) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_U45 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n281), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n267) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_U44 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n244), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n236), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n281) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_U43 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n235), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n234), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n233), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n242) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_U42 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n247), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n261), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n235), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n233) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_U41 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n266), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n232), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n231), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n234) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_U40 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n277), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n231) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_U39 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n257), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n237), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n277) );
  OR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_U38 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n268), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n238), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n237) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_U37 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n253), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n257) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_U36 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n239), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n268), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n232) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_U35 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n274), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n239) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_U34 ( .A(
        Red_StateRegOutput[28]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n230), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n287) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_U33 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n265), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n229), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n228), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n230) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_U32 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n247), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n249), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n227), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n226), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n228) );
  OR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_U31 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n235), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n261), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n255), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n226) );
  OR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_U30 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n274), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n238), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n248), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n255) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_U29 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n244), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n235) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_U28 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n253), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n236), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n252), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n225), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n238), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n227) );
  AND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_U27 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n253), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n236), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n225) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_U26 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n268), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n244), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n252) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_U25 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n251), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n274), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n236) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_U24 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n248), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n251) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_U23 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n265), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n266), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n253) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_U22 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n266), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n238), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n249) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_U21 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n261), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n266) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_U20 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n268), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n274), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n247) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_U19 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n245), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n268) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_U18 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n245), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n224), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n248), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n224), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n238), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n229) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_U17 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n223), .B(
        Red_StateRegOutput[28]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n238) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_U16 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n222), .B(
        F_SD2_RedSB_inst_n34), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n223) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_U15 ( .A(
        Red_StateRegOutput[30]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n222), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n248) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_U14 ( .A(
        F_SD2_RedSB_inst_n35), .B(F_SD2_RedSB_inst_n33), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n222) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_U13 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n244), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n274), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n261), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n224) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_U12 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n221), .B(
        Red_StateRegOutput[31]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n261) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_U11 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n220), .B(
        F_SD2_RedSB_inst_n34), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n274) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_U10 ( .A(
        Red_StateRegOutput[33]), .B(F_SD2_RedSB_inst_n36), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n220) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_U9 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n219), .B(
        Red_StateRegOutput[29]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n244) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_U8 ( .A(
        F_SD2_RedSB_inst_n34), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n221), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n219) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_U7 ( .A(
        F_SD2_RedSB_inst_n33), .B(F_SD2_RedSB_inst_n36), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n221) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_U6 ( .A(
        Red_StateRegOutput[34]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n218), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n245) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_U5 ( .A(
        F_SD2_RedSB_inst_n35), .B(F_SD2_RedSB_inst_n36), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n218) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_U4 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n217), .B(
        Red_StateRegOutput[32]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n265) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_U3 ( .A(
        F_SD2_RedSB_inst_n35), .B(F_SD2_RedSB_inst_n34), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_32_n217) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_U73 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n284), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n283), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n282), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n281), .ZN(Red_Feedback[61])
         );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_U72 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n280), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n281), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n279), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n283) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_U71 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n280), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n281), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n282), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n279) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_U70 ( .A(
        Red_StateRegOutput[33]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n278), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n282) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_U69 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n277), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n276), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n278) );
  NAND4_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_U68 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n275), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n274), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n273), .A4(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n272), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n276) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_U67 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n271), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n270), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n269), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n268), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n277) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_U66 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n267), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n268) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_U65 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n274), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n266), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n265), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n264), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n270) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_U64 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n263), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n265) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_U63 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n262), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n272), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n261), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n260), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n266) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_U62 ( .A(
        Red_StateRegOutput[29]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n259), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n281) );
  NOR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_U61 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n258), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n257), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n256), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n259) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_U60 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n255), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n254), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n255), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n253), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n252), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n256) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_U59 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n273), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n263), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n252) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_U58 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n251), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n250), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n263) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_U57 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n275), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n262), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n253) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_U56 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n271), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n269), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n254) );
  AOI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_U55 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n275), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n249), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n248), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n247), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n257) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_U54 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n246), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n245), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n275), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n247) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_U53 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n271), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n244), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n249) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_U52 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n245), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n271) );
  NOR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_U51 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n251), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n244), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n250), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n258) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_U50 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n260), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n248), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n250) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_U49 ( .A(
        Red_StateRegOutput[28]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n243), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n280) );
  AOI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_U48 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n275), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n242), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n241), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n240), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n243) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_U47 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n251), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n239), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n255), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n238), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n240) );
  OR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_U46 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n251), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n239), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n260), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n238) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_U45 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n237), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n248), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n244), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n255) );
  NOR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_U44 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n237), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n236), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n272), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n241) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_U43 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n274), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n262), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n246), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n235), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n236) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_U42 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n234), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n260), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n233), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n242) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_U41 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n232), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n246), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n262), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n233) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_U40 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n231), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n234) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_U39 ( .A(
        Red_StateRegOutput[30]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n230), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n284) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_U38 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n262), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n229), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n228), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n230) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_U37 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n267), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n227), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n226), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n264), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n228) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_U36 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n244), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n225), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n264) );
  NAND4_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_U35 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n237), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n269), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n274), .A4(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n227), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n226) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_U34 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n272), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n269) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_U33 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n237), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n273), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n262), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n231), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n267) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_U32 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n245), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n248), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n231) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_U31 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n244), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n239), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n273) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_U30 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n245), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n225), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n239) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_U29 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n260), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n237) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_U28 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n274), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n224), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n223), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n251), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n229) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_U27 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n232), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n244), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n261), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n244), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n235), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n224) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_U26 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n275), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n245), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n235) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_U25 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n227), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n275) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_U24 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n251), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n261) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_U23 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n227), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n272), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n251) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_U22 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n222), .B(
        Red_StateRegOutput[32]), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n272) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_U21 ( .A(
        F_SD2_RedSB_inst_n34), .B(F_SD2_RedSB_inst_n35), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n222) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_U20 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n221), .B(
        Red_StateRegOutput[31]), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n227) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_U19 ( .A(
        F_SD2_RedSB_inst_n33), .B(F_SD2_RedSB_inst_n36), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n221) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_U18 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n246), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n244) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_U17 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n220), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n219), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n246) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_U16 ( .A(
        F_SD2_RedSB_inst_n36), .B(Red_StateRegOutput[29]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n220) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_U15 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n223), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n232) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_U14 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n260), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n245), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n223) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_U13 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n218), .B(
        Red_StateRegOutput[33]), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n245) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_U12 ( .A(
        F_SD2_RedSB_inst_n34), .B(F_SD2_RedSB_inst_n36), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n218) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_U11 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n217), .B(
        F_SD2_RedSB_inst_n35), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n260) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_U10 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n219), .B(
        Red_StateRegOutput[28]), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n217) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_U9 ( .A(
        F_SD2_RedSB_inst_n33), .B(F_SD2_RedSB_inst_n34), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n219) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_U8 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n248), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n274) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_U7 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n216), .B(
        Red_StateRegOutput[34]), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n248) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_U6 ( .A(
        F_SD2_RedSB_inst_n35), .B(F_SD2_RedSB_inst_n36), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n216) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_U5 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n225), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n262) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_U4 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n215), .B(
        F_SD2_RedSB_inst_n35), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n225) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_U3 ( .A(
        Red_StateRegOutput[30]), .B(F_SD2_RedSB_inst_n33), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_33_n215) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_U65 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n283), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n282), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n281), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n280), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n279), .ZN(Red_Feedback[62])
         );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_U64 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n283), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n282), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n281), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n279) );
  MUX2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_U63 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n283), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n282), .S(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n278), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n280) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_U62 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n277), .B(
        Red_StateRegOutput[30]), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n278) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_U61 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n276), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n275), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n274), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n277) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_U60 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n273), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n274) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_U59 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n272), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n271), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n270), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n269), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n268), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n273) );
  AND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_U58 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n267), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n266), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n265), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n269) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_U57 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n266), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n264), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n263), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n262), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n275) );
  AOI222_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_U56 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n261), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n260), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n261), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n259), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n260), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n259), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n263) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_U55 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n258), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n268), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n259) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_U54 ( .A(
        Red_StateRegOutput[28]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n257), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n281) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_U53 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n268), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n256), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n255), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n257) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_U52 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n268), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n254), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n262), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n255) );
  AOI222_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_U51 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n261), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n260), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n261), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n253), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n260), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n253), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n254) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_U50 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n276), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n258), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n253) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_U49 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n252), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n251), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n250), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n249), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n256) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_U48 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n276), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n266), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n248), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n247), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n252) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_U47 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n264), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n247) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_U46 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n272), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n258), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n264) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_U45 ( .A(
        Red_StateRegOutput[29]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n246), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n282) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_U44 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n248), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n262), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n245), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n244), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n246) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_U43 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n248), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n243), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n244) );
  AOI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_U42 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n271), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n242), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n241), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n240), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n245) );
  NOR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_U41 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n270), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n239), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n250), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n240) );
  AND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_U40 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n238), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n268), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n260), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n241) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_U39 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n248), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n266), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n260) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_U38 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n251), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n237), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n249), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n238) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_U37 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n276), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n270), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n249) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_U36 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n258), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n236), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n262) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_U35 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n237), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n258) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_U34 ( .A(
        Red_StateRegOutput[33]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n235), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n283) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_U33 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n234), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n237), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n233), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n237), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n232), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n235) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_U32 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n251), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n268), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n267), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n236), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n271), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n232) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_U31 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n250), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n276), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n271) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_U30 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n237), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n248), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n250) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_U29 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n239), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n272), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n236) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_U28 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n242), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n265), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n243), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n233) );
  AND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_U27 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n261), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n231), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n243) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_U26 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n276), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n248), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n265) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_U25 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n230), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n229), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n248) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_U24 ( .A(
        F_SD2_RedSB_inst_n33), .B(Red_StateRegOutput[29]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n230) );
  OR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_U23 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n261), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n231), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n242) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_U22 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n268), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n266), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n231) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_U21 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n228), .B(
        Red_StateRegOutput[28]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n268) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_U20 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n227), .B(
        F_SD2_RedSB_inst_n34), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n228) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_U19 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n267), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n270), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n261) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_U18 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n272), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n270) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_U17 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n226), .B(
        Red_StateRegOutput[31]), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n272) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_U16 ( .A(
        F_SD2_RedSB_inst_n33), .B(F_SD2_RedSB_inst_n36), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n226) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_U15 ( .A(
        Red_StateRegOutput[33]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n229), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n237) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_U14 ( .A(
        F_SD2_RedSB_inst_n36), .B(F_SD2_RedSB_inst_n34), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n229) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_U13 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n225), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n234) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_U12 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n267), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n239), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n224), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n225) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_U11 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n267), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n239), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n276), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n224) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_U10 ( .A(
        Red_StateRegOutput[30]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n227), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n276) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_U9 ( .A(
        F_SD2_RedSB_inst_n35), .B(F_SD2_RedSB_inst_n33), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n227) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_U8 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n266), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n239) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_U7 ( .A(
        Red_StateRegOutput[34]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n223), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n266) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_U6 ( .A(
        F_SD2_RedSB_inst_n35), .B(F_SD2_RedSB_inst_n36), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n223) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_U5 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n251), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n267) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_U4 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n222), .B(
        Red_StateRegOutput[32]), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n251) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_U3 ( .A(
        F_SD2_RedSB_inst_n35), .B(F_SD2_RedSB_inst_n34), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_34_n222) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_U69 ( .A(
        Red_StateRegOutput[36]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n280), .Z(Red_Feedback[77])
         );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_U68 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n279), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n278), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n280) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_U67 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n277), .B2(
        Red_StateRegOutput[37]), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n276), .C2(
        Red_StateRegOutput[40]), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n275), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n278) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_U66 ( .A1(
        Red_StateRegOutput[37]), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n277), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n276), .B2(
        Red_StateRegOutput[40]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n275) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_U65 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n274), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n273), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n276) );
  AOI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_U64 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n272), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n271), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n270), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n269), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n273) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_U63 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n268), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n267), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n266), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n265), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n264), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n269) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_U62 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n268), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n263), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n262), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n270) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_U61 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n268), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n263), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n261), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n262) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_U60 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n260), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n259), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n258), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n271) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_U59 ( .A(
        Red_StateRegOutput[35]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n257), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n274) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_U58 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n253), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n254), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n251), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n255) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_U57 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n243), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n242), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n244), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n241), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n240), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n277) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_U56 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n239), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n238), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n237), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n240) );
  AOI222_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_U55 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n254), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n252), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n254), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n236), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n252), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n236), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n238) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_U54 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n246), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n267), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n236) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_U53 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n263), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n250), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n252) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_U52 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n235), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n254) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_U51 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n256), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n234), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n241) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_U50 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n261), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n263), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n233), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n242) );
  NOR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_U49 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n267), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n248), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n259), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n233) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_U48 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n249), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n250), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n259) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_U47 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n268), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n232), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n248) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_U46 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n256), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n267) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_U45 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n246), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n249), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n261) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_U44 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n264), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n260), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n231), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n279) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_U43 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n250), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n230), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n229), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n231) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_U42 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n250), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n228), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n251), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n229) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_U41 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n239), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n251) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_U40 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n246), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n265), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n239) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_U39 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n243), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n232), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n265) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_U38 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n245), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n247), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n256), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n263), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n228) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_U37 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n244), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n249), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n247) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_U36 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n266), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n246), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n245) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_U35 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n272), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n227), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n258), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n230) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_U34 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n235), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n226), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n258) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_U33 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n244), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n232), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n227) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_U32 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n235), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n226), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n260) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_U31 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n232), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n256), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n226) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_U30 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n225), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n224), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n256) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_U29 ( .A(
        Red_StateRegOutput[35]), .B(F_SD2_RedSB_inst_n37), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n225) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_U28 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n263), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n232) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_U27 ( .A(
        Red_StateRegOutput[41]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n223), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n263) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_U26 ( .A(
        F_SD2_RedSB_inst_n40), .B(F_SD2_RedSB_inst_n39), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n223) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_U25 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n243), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n268), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n235) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_U24 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n266), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n268) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_U23 ( .A(
        Red_StateRegOutput[39]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n224), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n266) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_U22 ( .A(
        F_SD2_RedSB_inst_n38), .B(F_SD2_RedSB_inst_n39), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n224) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_U21 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n244), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n243) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_U20 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n222), .B(
        Red_StateRegOutput[38]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n244) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_U19 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n234), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n264) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_U18 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n253), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n250), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n234) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_U17 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n221), .B(
        F_SD2_RedSB_inst_n38), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n250) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_U16 ( .A(
        Red_StateRegOutput[36]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n222), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n221) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_U15 ( .A(
        F_SD2_RedSB_inst_n40), .B(F_SD2_RedSB_inst_n37), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n222) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_U14 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n246), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n249), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n253) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_U13 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n237), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n249) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_U12 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n220), .B(
        Red_StateRegOutput[37]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n237) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_U11 ( .A(
        F_SD2_RedSB_inst_n37), .B(F_SD2_RedSB_inst_n39), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n220) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_U10 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n272), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n246) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_U9 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n219), .B(
        F_SD2_RedSB_inst_n38), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n272) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_U8 ( .A(
        Red_StateRegOutput[40]), .B(F_SD2_RedSB_inst_n40), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n219) );
  OAI33_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_U7 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n256), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n215), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n217), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n218), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n267), .B3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n255), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n257) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_U6 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n254), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n253), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n252), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n218) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_U5 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n250), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n216), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n217) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_U4 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n246), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n247), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n244), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n245), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n216) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_U3 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n249), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n248), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_35_n215) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_U68 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n273), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n274) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_U67 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n272), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n271), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n275) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_U66 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n267), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n266), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n269) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_U65 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n272), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n271), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n264), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n265) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_U64 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n260), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n259), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n267), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n268), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n261) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_U63 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n258), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n257), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n268) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_U62 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n256), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n267), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n255), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n254), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n260) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_U61 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n253), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n267) );
  NOR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_U60 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n252), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n251), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n250), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n262) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_U59 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n270), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n263) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_U58 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n258), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n257), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n270) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_U57 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n272), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n249), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n257) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_U56 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n252), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n273), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n246) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_U55 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n264), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n250), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n273) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_U54 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n253), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n259), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n250) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_U53 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n266), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n264) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_U52 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n252), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n259), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n248) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_U51 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n278), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n259) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_U50 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n278), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n249), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n245) );
  AND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_U49 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n277), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n271), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n258) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_U48 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n272), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n253), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n255) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_U47 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n251), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n272) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_U46 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n251), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n277), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n256) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_U45 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n252), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n277) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_U44 ( .A(
        Red_StateRegOutput[40]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n244), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n278) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_U43 ( .A(
        F_SD2_RedSB_inst_n39), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n243), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n266) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_U42 ( .A(
        Red_StateRegOutput[37]), .B(F_SD2_RedSB_inst_n37), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n243) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_U41 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n254), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n276) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_U40 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n271), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n247), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n254) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_U39 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n249), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n247) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_U38 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n242), .B(
        Red_StateRegOutput[35]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n249) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_U37 ( .A(
        F_SD2_RedSB_inst_n37), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n241), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n242) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_U36 ( .A(
        Red_StateRegOutput[39]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n241), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n271) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_U35 ( .A(
        F_SD2_RedSB_inst_n39), .B(F_SD2_RedSB_inst_n38), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n241) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_U34 ( .A(
        Red_StateRegOutput[41]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n240), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n251) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_U33 ( .A(
        F_SD2_RedSB_inst_n39), .B(F_SD2_RedSB_inst_n40), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n240) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_U32 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n239), .B(
        Red_StateRegOutput[38]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n252) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_U31 ( .A(
        F_SD2_RedSB_inst_n37), .B(F_SD2_RedSB_inst_n40), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n239) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_U30 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n238), .B(
        Red_StateRegOutput[36]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n253) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_U29 ( .A(
        F_SD2_RedSB_inst_n37), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n244), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n238) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_U28 ( .A(
        F_SD2_RedSB_inst_n38), .B(F_SD2_RedSB_inst_n40), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n244) );
  AOI222_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_U27 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n221), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n228), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n221), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n233), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n228), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n237), .ZN(Red_Feedback[78])
         );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_U26 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n236), .B(
        Red_StateRegOutput[36]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n237) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_U25 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n234), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n235), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n236) );
  AOI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_U24 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n273), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n263), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n261), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n262), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n235) );
  NAND4_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_U23 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n249), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n252), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n264), .A4(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n255), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n234) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_U22 ( .A(
        Red_StateRegOutput[40]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n232), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n233) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_U21 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n229), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n278), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n230), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n278), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n231), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n232) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_U20 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n277), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n276), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n275), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n276), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n274), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n231) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_U19 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n270), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n269), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n268), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n230) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_U18 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n272), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n271), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n265), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n229) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_U17 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n227), .B(
        Red_StateRegOutput[37]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n228) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_U16 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n266), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n222), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n226), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n227) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_U15 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n247), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n246), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n225), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n226) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_U14 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n224), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n255), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n224), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n245), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n264), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n225) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_U13 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n217), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n223), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n224) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_U12 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n251), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n248), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n258), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n245), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n223) );
  NOR4_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_U11 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n251), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n252), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n253), .A4(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n276), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n222) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_U10 ( .A(
        Red_StateRegOutput[35]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n220), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n221) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_U9 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n249), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n216), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n219), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n220) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_U8 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n249), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n217), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n218), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n219) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_U7 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n258), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n255), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n259), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n266), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n218) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_U6 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n278), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n256), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n258), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n255), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n217) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_U5 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n250), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n214), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n271), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n215), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n216) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_U4 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n264), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n272), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n253), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n248), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n215) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_U3 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n252), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n264), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_36_n214) );
  MUX2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_U54 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n240), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n239), .S(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n238), .Z(Red_Feedback[79])
         );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_U53 ( .A(
        Red_StateRegOutput[37]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n237), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n238) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_U52 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n236), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n235), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n234), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n233), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n237) );
  OR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_U51 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n232), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n231), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n230), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n233) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_U50 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n229), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n228), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n227), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n234) );
  AOI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_U49 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n226), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n225), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n224), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n223), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n236) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_U48 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n222), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n221), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n220), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n221), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n219), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n223) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_U47 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n226), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n225), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n218), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n221) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_U46 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n217), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n216), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n225) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_U45 ( .A(
        Red_StateRegOutput[40]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n215), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n239) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_U44 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n214), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n230), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n213), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n212), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n215) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_U43 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n228), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n226), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n211), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n232), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n212) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_U42 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n210), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n228), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n210), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n226), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n216), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n213) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_U41 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n220), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n216) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_U40 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n209), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n226) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_U39 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n208), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n207), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n228) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_U38 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n219), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n206), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n205), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n210) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_U37 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n219), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n206), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n208), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n205) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_U36 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n235), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n208) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_U35 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n222), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n204), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n229), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n214) );
  AND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_U34 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n206), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n219), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n204) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_U33 ( .A(
        Red_StateRegOutput[36]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n203), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n240) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_U32 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n202), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n201), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n200), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n201), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n199), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n203) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_U31 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n198), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n197), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n230), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n209), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n199) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_U30 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n227), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n220), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n218), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n197) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_U29 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n207), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n218) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_U28 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n222), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n201), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n227) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_U27 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n198), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n230), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n209), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n230), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n217), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n200) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_U26 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n231), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n206), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n209) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_U25 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n207), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n235), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n220), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n230) );
  AOI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_U24 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n229), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n211), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n207), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n224), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n198) );
  NOR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_U23 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n231), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n220), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n201), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n224) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_U22 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n219), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n220), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n211) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_U21 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n196), .B(
        Red_StateRegOutput[40]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n220) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_U20 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n201), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n219) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_U19 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n232), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n206), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n229) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_U18 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n195), .B(
        Red_StateRegOutput[39]), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n206) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_U17 ( .A(
        F_SD2_RedSB_inst_n39), .B(F_SD2_RedSB_inst_n38), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n195) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_U16 ( .A(
        Red_StateRegOutput[41]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n194), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n201) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_U15 ( .A(
        F_SD2_RedSB_inst_n39), .B(F_SD2_RedSB_inst_n40), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n194) );
  NOR4_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_U14 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n207), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n231), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n232), .A4(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n235), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n202) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_U13 ( .A(
        Red_StateRegOutput[37]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n193), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n235) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_U12 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n217), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n232) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_U11 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n192), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n193), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n217) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_U10 ( .A(
        F_SD2_RedSB_inst_n37), .B(F_SD2_RedSB_inst_n39), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n193) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_U9 ( .A(
        F_SD2_RedSB_inst_n38), .B(Red_StateRegOutput[35]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n192) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_U8 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n222), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n231) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_U7 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n191), .B(
        Red_StateRegOutput[38]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n222) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_U6 ( .A(
        F_SD2_RedSB_inst_n37), .B(F_SD2_RedSB_inst_n40), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n191) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_U5 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n190), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n196), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n207) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_U4 ( .A(
        F_SD2_RedSB_inst_n38), .B(F_SD2_RedSB_inst_n40), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n196) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_U3 ( .A(
        F_SD2_RedSB_inst_n37), .B(Red_StateRegOutput[36]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_37_n190) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_U69 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n289), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n288), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n287), .ZN(Red_Feedback[80])
         );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_U68 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n285), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n284), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n283), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n288) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_U67 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n284), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n286), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n285), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n283) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_U66 ( .A(
        Red_StateRegOutput[40]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n270), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n284) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_U65 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n269), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n268), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n267), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n271), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n270) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_U64 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n266), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n276), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n265), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n264), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n263), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n267) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_U63 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n262), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n261), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n280), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n260), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n265) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_U62 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n264), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n276) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_U61 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n275), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n274), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n266) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_U60 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n259), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n268) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_U59 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n258), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n257), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n256), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n269) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_U58 ( .A(
        Red_StateRegOutput[37]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n255), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n285) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_U57 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n254), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n264), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n253), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n252), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n255) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_U56 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n280), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n259), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n251), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n252) );
  NAND4_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_U55 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n256), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n250), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n278), .A4(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n264), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n253) );
  AOI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_U54 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n273), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n249), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n248), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n279), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n254) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_U53 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n260), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n261), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n247), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n279) );
  NOR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_U52 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n280), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n246), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n282), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n248) );
  AND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_U51 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n260), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n261), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n282) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_U50 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n245), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n261) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_U49 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n251), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n271), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n273) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_U48 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n278), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n281), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n259) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_U47 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n264), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n271), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n281) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_U46 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n246), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n258), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n247) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_U45 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n243), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n249), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n258) );
  AND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_U44 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n245), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n244), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n263) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_U43 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n280), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n274), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n244) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_U42 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n251), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n275), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n245) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_U41 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n257), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n275) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_U40 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n251), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n249), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n250) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_U39 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n277), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n257), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n256) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_U38 ( .A(
        Red_StateRegOutput[39]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n242), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n257) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_U37 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n280), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n277) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_U36 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n271), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n246) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_U35 ( .A(
        Red_StateRegOutput[40]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n241), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n271) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_U34 ( .A(
        F_SD2_RedSB_inst_n38), .B(F_SD2_RedSB_inst_n40), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n241) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_U33 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n264), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n243), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n272) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_U32 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n251), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n243) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_U31 ( .A(
        Red_StateRegOutput[38]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n240), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n251) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_U30 ( .A(
        F_SD2_RedSB_inst_n37), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n239), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n264) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_U29 ( .A(
        Red_StateRegOutput[37]), .B(F_SD2_RedSB_inst_n39), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n239) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_U28 ( .A(
        F_SD2_RedSB_inst_n38), .B(F_SD2_RedSB_inst_n39), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n242) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_U27 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n278), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n249), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n260) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_U26 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n274), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n249) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_U25 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n238), .B(
        Red_StateRegOutput[41]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n274) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_U24 ( .A(
        F_SD2_RedSB_inst_n39), .B(F_SD2_RedSB_inst_n40), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n238) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_U23 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n262), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n278) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_U22 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n237), .B(
        Red_StateRegOutput[36]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n262) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_U21 ( .A(
        F_SD2_RedSB_inst_n38), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n240), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n237) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_U20 ( .A(
        F_SD2_RedSB_inst_n37), .B(F_SD2_RedSB_inst_n40), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n240) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_U19 ( .A(
        Red_StateRegOutput[36]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n236), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n289) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_U18 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n260), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n232), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n234), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n235), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n236) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_U17 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n263), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n271), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n263), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n250), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n262), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n235) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_U16 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n245), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n259), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n244), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n259), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n233), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n234) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_U15 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n262), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n247), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n233) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_U14 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n280), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n272), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n246), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n256), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n232) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_U13 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n286), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n288), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n230), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n231), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n289), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n287) );
  OR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_U12 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n285), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n284), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n231) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_U11 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n286), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n230) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_U10 ( .A(
        Red_StateRegOutput[35]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n229), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n280) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_U9 ( .A(
        F_SD2_RedSB_inst_n37), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n242), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n229) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_U8 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n228), .B(
        Red_StateRegOutput[35]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n286) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_U7 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n224), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n279), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n227), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n228) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_U6 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n278), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n225), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n277), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n226), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n227) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_U5 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n276), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n274), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n275), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n226) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_U4 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n271), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n272), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n275), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n273), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n225) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_U3 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n282), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n281), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n280), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_38_n224) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_U73 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n277), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n276), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n279), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n278) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_U72 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n275), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n274), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n273), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n277) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_U71 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n272), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n279) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_U70 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n266), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n265), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n264), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n267) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_U69 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n265), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n269) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_U68 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n280), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n263) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_U67 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n261), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n260), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n280) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_U66 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n264), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n281), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n258), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n276) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_U65 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n283), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n275), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n259) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_U64 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n264), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n257), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n283) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_U63 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n261), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n262), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n254), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n285), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n255) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_U62 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n272), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n253), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n285) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_U61 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n270), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n252), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n282) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_U60 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n286), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n274) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_U59 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n257), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n251), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n286) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_U58 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n250), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n249), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n248), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n256) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_U57 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n260), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n271), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n250), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n248) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_U56 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n273), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n247), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n246), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n249) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_U55 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n284), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n246) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_U54 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n270), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n252), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n284) );
  OR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_U53 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n275), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n253), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n252) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_U52 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n266), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n270) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_U51 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n254), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n275), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n247) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_U50 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n281), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n254) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_U49 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n272), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n244), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n243), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n245) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_U48 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n260), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n262), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n242), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n241), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n243) );
  OR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_U47 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n250), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n271), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n268), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n241) );
  OR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_U46 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n281), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n253), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n261), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n268) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_U45 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n257), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n250) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_U44 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n266), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n251), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n265), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n240), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n253), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n242) );
  AND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_U43 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n266), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n251), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n240) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_U42 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n275), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n257), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n265) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_U41 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n264), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n281), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n251) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_U40 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n261), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n264) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_U39 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n272), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n273), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n266) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_U38 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n273), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n253), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n262) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_U37 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n271), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n273) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_U36 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n275), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n281), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n260) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_U35 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n258), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n275) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_U34 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n258), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n239), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n261), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n239), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n253), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n244) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_U33 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n238), .B(
        Red_StateRegOutput[35]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n253) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_U32 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n237), .B(
        F_SD2_RedSB_inst_n38), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n238) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_U31 ( .A(
        Red_StateRegOutput[37]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n237), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n261) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_U30 ( .A(
        F_SD2_RedSB_inst_n39), .B(F_SD2_RedSB_inst_n37), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n237) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_U29 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n257), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n281), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n271), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n239) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_U28 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n236), .B(
        Red_StateRegOutput[38]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n271) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_U27 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n235), .B(
        F_SD2_RedSB_inst_n38), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n281) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_U26 ( .A(
        Red_StateRegOutput[40]), .B(F_SD2_RedSB_inst_n40), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n235) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_U25 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n234), .B(
        Red_StateRegOutput[36]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n257) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_U24 ( .A(
        F_SD2_RedSB_inst_n38), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n236), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n234) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_U23 ( .A(
        F_SD2_RedSB_inst_n37), .B(F_SD2_RedSB_inst_n40), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n236) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_U22 ( .A(
        Red_StateRegOutput[41]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n233), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n258) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_U21 ( .A(
        F_SD2_RedSB_inst_n39), .B(F_SD2_RedSB_inst_n40), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n233) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_U20 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n232), .B(
        Red_StateRegOutput[39]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n272) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_U19 ( .A(
        F_SD2_RedSB_inst_n39), .B(F_SD2_RedSB_inst_n38), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n232) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_U18 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n217), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n220), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n230), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n224), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n231), .ZN(Red_Feedback[81])
         );
  NOR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_U17 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n220), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n224), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n230), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n231) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_U16 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n228), .B2(
        Red_StateRegOutput[37]), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n229), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n230) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_U15 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n228), .B2(
        Red_StateRegOutput[37]), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n217), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n229) );
  AOI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_U14 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n271), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n225), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n226), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n227), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n228) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_U13 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n262), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n286), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n263), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n271), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n227) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_U12 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n270), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n269), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n267), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n268), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n226) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_U11 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n285), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n259), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n276), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n225) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_U10 ( .A(
        Red_StateRegOutput[40]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n223), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n224) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_U9 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n285), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n286), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n221), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n222), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n223) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_U8 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n279), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n280), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n278), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n222) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_U7 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n284), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n282), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n284), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n283), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n281), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n221) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_U6 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n219), .B(
        Red_StateRegOutput[36]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n220) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_U5 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n218), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n256), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n219) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_U4 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n265), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n255), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n282), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n274), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n218) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_U3 ( .A(
        Red_StateRegOutput[35]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n245), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_39_n217) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_U73 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n284), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n283), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n282), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n281), .ZN(Red_Feedback[82])
         );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_U72 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n280), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n281), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n279), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n283) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_U71 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n280), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n281), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n282), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n279) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_U70 ( .A(
        Red_StateRegOutput[40]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n278), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n282) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_U69 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n277), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n276), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n278) );
  NAND4_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_U68 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n275), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n274), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n273), .A4(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n272), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n276) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_U67 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n271), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n270), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n269), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n268), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n277) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_U66 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n267), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n268) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_U65 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n274), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n266), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n265), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n264), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n270) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_U64 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n263), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n265) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_U63 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n262), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n272), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n261), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n260), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n266) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_U62 ( .A(
        Red_StateRegOutput[36]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n259), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n281) );
  NOR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_U61 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n258), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n257), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n256), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n259) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_U60 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n255), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n254), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n255), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n253), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n252), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n256) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_U59 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n273), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n263), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n252) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_U58 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n251), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n250), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n263) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_U57 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n275), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n262), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n253) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_U56 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n271), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n269), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n254) );
  AOI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_U55 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n275), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n249), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n248), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n247), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n257) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_U54 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n246), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n245), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n275), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n247) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_U53 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n271), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n244), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n249) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_U52 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n245), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n271) );
  NOR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_U51 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n251), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n244), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n250), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n258) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_U50 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n260), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n248), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n250) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_U49 ( .A(
        Red_StateRegOutput[35]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n243), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n280) );
  AOI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_U48 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n275), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n242), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n241), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n240), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n243) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_U47 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n251), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n239), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n255), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n238), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n240) );
  OR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_U46 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n251), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n239), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n260), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n238) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_U45 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n237), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n248), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n244), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n255) );
  NOR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_U44 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n237), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n236), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n272), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n241) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_U43 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n274), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n262), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n246), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n235), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n236) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_U42 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n234), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n260), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n233), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n242) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_U41 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n232), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n246), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n262), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n233) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_U40 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n231), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n234) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_U39 ( .A(
        Red_StateRegOutput[37]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n230), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n284) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_U38 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n262), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n229), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n228), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n230) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_U37 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n267), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n227), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n226), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n264), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n228) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_U36 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n244), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n225), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n264) );
  NAND4_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_U35 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n237), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n269), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n274), .A4(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n227), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n226) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_U34 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n272), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n269) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_U33 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n237), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n273), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n262), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n231), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n267) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_U32 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n245), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n248), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n231) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_U31 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n244), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n239), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n273) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_U30 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n245), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n225), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n239) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_U29 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n260), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n237) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_U28 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n274), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n224), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n223), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n251), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n229) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_U27 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n232), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n244), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n261), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n244), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n235), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n224) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_U26 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n275), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n245), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n235) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_U25 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n227), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n275) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_U24 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n251), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n261) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_U23 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n227), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n272), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n251) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_U22 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n222), .B(
        Red_StateRegOutput[39]), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n272) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_U21 ( .A(
        F_SD2_RedSB_inst_n38), .B(F_SD2_RedSB_inst_n39), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n222) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_U20 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n221), .B(
        Red_StateRegOutput[38]), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n227) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_U19 ( .A(
        F_SD2_RedSB_inst_n37), .B(F_SD2_RedSB_inst_n40), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n221) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_U18 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n246), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n244) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_U17 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n220), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n219), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n246) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_U16 ( .A(
        F_SD2_RedSB_inst_n40), .B(Red_StateRegOutput[36]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n220) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_U15 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n223), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n232) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_U14 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n260), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n245), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n223) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_U13 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n218), .B(
        Red_StateRegOutput[40]), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n245) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_U12 ( .A(
        F_SD2_RedSB_inst_n38), .B(F_SD2_RedSB_inst_n40), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n218) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_U11 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n217), .B(
        F_SD2_RedSB_inst_n39), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n260) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_U10 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n219), .B(
        Red_StateRegOutput[35]), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n217) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_U9 ( .A(
        F_SD2_RedSB_inst_n37), .B(F_SD2_RedSB_inst_n38), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n219) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_U8 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n248), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n274) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_U7 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n216), .B(
        Red_StateRegOutput[41]), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n248) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_U6 ( .A(
        F_SD2_RedSB_inst_n39), .B(F_SD2_RedSB_inst_n40), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n216) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_U5 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n225), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n262) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_U4 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n215), .B(
        F_SD2_RedSB_inst_n39), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n225) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_U3 ( .A(
        Red_StateRegOutput[37]), .B(F_SD2_RedSB_inst_n37), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_40_n215) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_U65 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n283), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n282), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n281), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n280), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n279), .ZN(Red_Feedback[83])
         );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_U64 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n283), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n282), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n281), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n279) );
  MUX2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_U63 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n283), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n282), .S(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n278), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n280) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_U62 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n277), .B(
        Red_StateRegOutput[37]), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n278) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_U61 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n276), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n275), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n274), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n277) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_U60 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n273), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n274) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_U59 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n272), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n271), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n270), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n269), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n268), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n273) );
  AND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_U58 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n267), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n266), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n265), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n269) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_U57 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n266), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n264), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n263), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n262), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n275) );
  AOI222_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_U56 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n261), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n260), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n261), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n259), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n260), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n259), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n263) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_U55 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n258), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n268), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n259) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_U54 ( .A(
        Red_StateRegOutput[35]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n257), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n281) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_U53 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n268), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n256), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n255), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n257) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_U52 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n268), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n254), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n262), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n255) );
  AOI222_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_U51 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n261), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n260), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n261), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n253), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n260), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n253), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n254) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_U50 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n276), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n258), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n253) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_U49 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n252), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n251), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n250), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n249), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n256) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_U48 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n276), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n266), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n248), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n247), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n252) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_U47 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n264), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n247) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_U46 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n272), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n258), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n264) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_U45 ( .A(
        Red_StateRegOutput[36]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n246), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n282) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_U44 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n248), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n262), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n245), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n244), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n246) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_U43 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n248), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n243), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n244) );
  AOI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_U42 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n271), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n242), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n241), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n240), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n245) );
  NOR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_U41 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n270), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n239), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n250), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n240) );
  AND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_U40 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n238), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n268), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n260), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n241) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_U39 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n248), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n266), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n260) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_U38 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n251), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n237), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n249), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n238) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_U37 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n276), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n270), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n249) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_U36 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n258), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n236), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n262) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_U35 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n237), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n258) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_U34 ( .A(
        Red_StateRegOutput[40]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n235), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n283) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_U33 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n234), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n237), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n233), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n237), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n232), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n235) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_U32 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n251), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n268), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n267), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n236), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n271), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n232) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_U31 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n250), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n276), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n271) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_U30 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n237), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n248), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n250) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_U29 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n239), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n272), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n236) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_U28 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n242), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n265), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n243), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n233) );
  AND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_U27 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n261), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n231), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n243) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_U26 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n276), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n248), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n265) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_U25 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n230), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n229), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n248) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_U24 ( .A(
        F_SD2_RedSB_inst_n37), .B(Red_StateRegOutput[36]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n230) );
  OR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_U23 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n261), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n231), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n242) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_U22 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n268), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n266), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n231) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_U21 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n228), .B(
        Red_StateRegOutput[35]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n268) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_U20 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n227), .B(
        F_SD2_RedSB_inst_n38), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n228) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_U19 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n267), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n270), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n261) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_U18 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n272), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n270) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_U17 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n226), .B(
        Red_StateRegOutput[38]), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n272) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_U16 ( .A(
        F_SD2_RedSB_inst_n37), .B(F_SD2_RedSB_inst_n40), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n226) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_U15 ( .A(
        Red_StateRegOutput[40]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n229), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n237) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_U14 ( .A(
        F_SD2_RedSB_inst_n40), .B(F_SD2_RedSB_inst_n38), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n229) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_U13 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n225), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n234) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_U12 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n267), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n239), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n224), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n225) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_U11 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n267), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n239), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n276), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n224) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_U10 ( .A(
        Red_StateRegOutput[37]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n227), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n276) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_U9 ( .A(
        F_SD2_RedSB_inst_n39), .B(F_SD2_RedSB_inst_n37), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n227) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_U8 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n266), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n239) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_U7 ( .A(
        Red_StateRegOutput[41]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n223), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n266) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_U6 ( .A(
        F_SD2_RedSB_inst_n39), .B(F_SD2_RedSB_inst_n40), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n223) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_U5 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n251), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n267) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_U4 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n222), .B(
        Red_StateRegOutput[39]), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n251) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_U3 ( .A(
        F_SD2_RedSB_inst_n39), .B(F_SD2_RedSB_inst_n38), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_41_n222) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_U69 ( .A(
        Red_StateRegOutput[43]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n280), .Z(Red_Feedback[70])
         );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_U68 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n279), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n278), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n280) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_U67 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n277), .B2(
        Red_StateRegOutput[44]), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n276), .C2(
        Red_StateRegOutput[47]), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n275), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n278) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_U66 ( .A1(
        Red_StateRegOutput[44]), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n277), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n276), .B2(
        Red_StateRegOutput[47]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n275) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_U65 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n274), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n273), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n276) );
  AOI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_U64 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n272), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n271), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n270), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n269), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n273) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_U63 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n268), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n267), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n266), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n265), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n264), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n269) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_U62 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n268), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n263), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n262), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n270) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_U61 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n268), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n263), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n261), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n262) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_U60 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n260), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n259), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n258), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n271) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_U59 ( .A(
        Red_StateRegOutput[42]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n257), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n274) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_U58 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n253), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n254), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n251), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n255) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_U57 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n243), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n242), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n244), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n241), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n240), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n277) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_U56 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n239), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n238), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n237), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n240) );
  AOI222_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_U55 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n254), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n252), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n254), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n236), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n252), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n236), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n238) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_U54 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n246), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n267), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n236) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_U53 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n263), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n250), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n252) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_U52 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n235), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n254) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_U51 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n256), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n234), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n241) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_U50 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n261), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n263), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n233), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n242) );
  NOR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_U49 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n267), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n248), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n259), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n233) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_U48 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n249), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n250), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n259) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_U47 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n268), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n232), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n248) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_U46 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n256), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n267) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_U45 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n246), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n249), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n261) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_U44 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n264), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n260), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n231), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n279) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_U43 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n250), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n230), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n229), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n231) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_U42 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n250), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n228), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n251), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n229) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_U41 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n239), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n251) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_U40 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n246), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n265), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n239) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_U39 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n243), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n232), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n265) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_U38 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n245), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n247), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n256), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n263), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n228) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_U37 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n244), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n249), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n247) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_U36 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n266), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n246), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n245) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_U35 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n272), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n227), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n258), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n230) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_U34 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n235), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n226), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n258) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_U33 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n244), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n232), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n227) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_U32 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n235), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n226), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n260) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_U31 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n232), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n256), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n226) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_U30 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n225), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n224), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n256) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_U29 ( .A(
        Red_StateRegOutput[42]), .B(F_SD2_RedSB_inst_n41), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n225) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_U28 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n263), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n232) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_U27 ( .A(
        Red_StateRegOutput[48]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n223), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n263) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_U26 ( .A(
        F_SD2_RedSB_inst_n44), .B(F_SD2_RedSB_inst_n43), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n223) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_U25 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n243), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n268), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n235) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_U24 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n266), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n268) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_U23 ( .A(
        Red_StateRegOutput[46]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n224), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n266) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_U22 ( .A(
        F_SD2_RedSB_inst_n42), .B(F_SD2_RedSB_inst_n43), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n224) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_U21 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n244), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n243) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_U20 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n222), .B(
        Red_StateRegOutput[45]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n244) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_U19 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n234), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n264) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_U18 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n253), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n250), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n234) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_U17 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n221), .B(
        F_SD2_RedSB_inst_n42), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n250) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_U16 ( .A(
        Red_StateRegOutput[43]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n222), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n221) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_U15 ( .A(
        F_SD2_RedSB_inst_n44), .B(F_SD2_RedSB_inst_n41), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n222) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_U14 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n246), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n249), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n253) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_U13 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n237), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n249) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_U12 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n220), .B(
        Red_StateRegOutput[44]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n237) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_U11 ( .A(
        F_SD2_RedSB_inst_n41), .B(F_SD2_RedSB_inst_n43), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n220) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_U10 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n272), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n246) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_U9 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n219), .B(
        F_SD2_RedSB_inst_n42), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n272) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_U8 ( .A(
        Red_StateRegOutput[47]), .B(F_SD2_RedSB_inst_n44), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n219) );
  OAI33_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_U7 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n256), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n215), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n217), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n218), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n267), .B3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n255), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n257) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_U6 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n254), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n253), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n252), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n218) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_U5 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n250), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n216), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n217) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_U4 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n246), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n247), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n244), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n245), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n216) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_U3 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n249), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n248), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_42_n215) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_U68 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n273), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n274) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_U67 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n272), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n271), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n275) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_U66 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n267), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n266), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n269) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_U65 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n272), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n271), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n264), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n265) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_U64 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n260), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n259), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n267), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n268), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n261) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_U63 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n258), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n257), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n268) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_U62 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n256), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n267), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n255), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n254), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n260) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_U61 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n253), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n267) );
  NOR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_U60 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n252), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n251), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n250), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n262) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_U59 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n270), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n263) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_U58 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n258), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n257), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n270) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_U57 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n272), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n249), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n257) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_U56 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n252), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n273), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n246) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_U55 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n264), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n250), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n273) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_U54 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n253), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n259), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n250) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_U53 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n266), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n264) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_U52 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n252), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n259), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n248) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_U51 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n278), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n259) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_U50 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n278), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n249), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n245) );
  AND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_U49 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n277), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n271), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n258) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_U48 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n272), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n253), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n255) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_U47 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n251), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n272) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_U46 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n251), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n277), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n256) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_U45 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n252), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n277) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_U44 ( .A(
        Red_StateRegOutput[47]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n244), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n278) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_U43 ( .A(
        F_SD2_RedSB_inst_n43), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n243), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n266) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_U42 ( .A(
        Red_StateRegOutput[44]), .B(F_SD2_RedSB_inst_n41), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n243) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_U41 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n254), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n276) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_U40 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n271), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n247), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n254) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_U39 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n249), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n247) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_U38 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n242), .B(
        Red_StateRegOutput[42]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n249) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_U37 ( .A(
        F_SD2_RedSB_inst_n41), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n241), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n242) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_U36 ( .A(
        Red_StateRegOutput[46]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n241), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n271) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_U35 ( .A(
        F_SD2_RedSB_inst_n43), .B(F_SD2_RedSB_inst_n42), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n241) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_U34 ( .A(
        Red_StateRegOutput[48]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n240), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n251) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_U33 ( .A(
        F_SD2_RedSB_inst_n43), .B(F_SD2_RedSB_inst_n44), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n240) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_U32 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n239), .B(
        Red_StateRegOutput[45]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n252) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_U31 ( .A(
        F_SD2_RedSB_inst_n41), .B(F_SD2_RedSB_inst_n44), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n239) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_U30 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n238), .B(
        Red_StateRegOutput[43]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n253) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_U29 ( .A(
        F_SD2_RedSB_inst_n41), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n244), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n238) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_U28 ( .A(
        F_SD2_RedSB_inst_n42), .B(F_SD2_RedSB_inst_n44), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n244) );
  AOI222_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_U27 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n221), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n228), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n221), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n233), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n228), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n237), .ZN(Red_Feedback[71])
         );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_U26 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n236), .B(
        Red_StateRegOutput[43]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n237) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_U25 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n234), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n235), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n236) );
  AOI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_U24 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n273), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n263), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n261), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n262), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n235) );
  NAND4_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_U23 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n249), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n252), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n264), .A4(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n255), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n234) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_U22 ( .A(
        Red_StateRegOutput[47]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n232), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n233) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_U21 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n229), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n278), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n230), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n278), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n231), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n232) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_U20 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n277), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n276), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n275), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n276), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n274), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n231) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_U19 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n270), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n269), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n268), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n230) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_U18 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n272), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n271), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n265), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n229) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_U17 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n227), .B(
        Red_StateRegOutput[44]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n228) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_U16 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n266), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n222), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n226), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n227) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_U15 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n247), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n246), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n225), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n226) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_U14 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n224), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n255), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n224), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n245), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n264), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n225) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_U13 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n217), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n223), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n224) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_U12 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n251), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n248), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n258), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n245), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n223) );
  NOR4_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_U11 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n251), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n252), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n253), .A4(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n276), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n222) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_U10 ( .A(
        Red_StateRegOutput[42]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n220), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n221) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_U9 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n249), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n216), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n219), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n220) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_U8 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n249), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n217), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n218), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n219) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_U7 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n258), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n255), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n259), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n266), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n218) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_U6 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n278), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n256), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n258), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n255), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n217) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_U5 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n250), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n214), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n271), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n215), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n216) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_U4 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n264), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n272), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n253), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n248), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n215) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_U3 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n252), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n264), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_43_n214) );
  MUX2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_U54 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n240), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n239), .S(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n238), .Z(Red_Feedback[72])
         );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_U53 ( .A(
        Red_StateRegOutput[44]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n237), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n238) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_U52 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n236), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n235), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n234), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n233), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n237) );
  OR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_U51 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n232), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n231), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n230), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n233) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_U50 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n229), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n228), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n227), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n234) );
  AOI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_U49 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n226), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n225), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n224), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n223), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n236) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_U48 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n222), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n221), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n220), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n221), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n219), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n223) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_U47 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n226), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n225), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n218), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n221) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_U46 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n217), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n216), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n225) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_U45 ( .A(
        Red_StateRegOutput[47]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n215), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n239) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_U44 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n214), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n230), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n213), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n212), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n215) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_U43 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n228), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n226), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n211), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n232), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n212) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_U42 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n210), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n228), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n210), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n226), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n216), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n213) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_U41 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n220), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n216) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_U40 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n209), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n226) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_U39 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n208), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n207), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n228) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_U38 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n219), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n206), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n205), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n210) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_U37 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n219), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n206), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n208), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n205) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_U36 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n235), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n208) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_U35 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n222), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n204), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n229), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n214) );
  AND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_U34 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n206), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n219), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n204) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_U33 ( .A(
        Red_StateRegOutput[43]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n203), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n240) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_U32 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n202), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n201), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n200), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n201), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n199), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n203) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_U31 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n198), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n197), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n230), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n209), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n199) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_U30 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n227), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n220), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n218), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n197) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_U29 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n207), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n218) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_U28 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n222), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n201), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n227) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_U27 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n198), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n230), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n209), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n230), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n217), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n200) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_U26 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n231), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n206), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n209) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_U25 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n207), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n235), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n220), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n230) );
  AOI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_U24 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n229), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n211), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n207), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n224), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n198) );
  NOR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_U23 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n231), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n220), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n201), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n224) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_U22 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n219), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n220), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n211) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_U21 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n196), .B(
        Red_StateRegOutput[47]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n220) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_U20 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n201), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n219) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_U19 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n232), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n206), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n229) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_U18 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n195), .B(
        Red_StateRegOutput[46]), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n206) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_U17 ( .A(
        F_SD2_RedSB_inst_n43), .B(F_SD2_RedSB_inst_n42), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n195) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_U16 ( .A(
        Red_StateRegOutput[48]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n194), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n201) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_U15 ( .A(
        F_SD2_RedSB_inst_n43), .B(F_SD2_RedSB_inst_n44), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n194) );
  NOR4_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_U14 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n207), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n231), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n232), .A4(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n235), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n202) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_U13 ( .A(
        Red_StateRegOutput[44]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n193), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n235) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_U12 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n217), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n232) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_U11 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n192), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n193), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n217) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_U10 ( .A(
        F_SD2_RedSB_inst_n41), .B(F_SD2_RedSB_inst_n43), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n193) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_U9 ( .A(
        F_SD2_RedSB_inst_n42), .B(Red_StateRegOutput[42]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n192) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_U8 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n222), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n231) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_U7 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n191), .B(
        Red_StateRegOutput[45]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n222) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_U6 ( .A(
        F_SD2_RedSB_inst_n41), .B(F_SD2_RedSB_inst_n44), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n191) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_U5 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n190), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n196), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n207) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_U4 ( .A(
        F_SD2_RedSB_inst_n42), .B(F_SD2_RedSB_inst_n44), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n196) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_U3 ( .A(
        F_SD2_RedSB_inst_n41), .B(Red_StateRegOutput[43]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_44_n190) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_U69 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n289), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n288), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n287), .ZN(Red_Feedback[73])
         );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_U68 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n285), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n284), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n283), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n288) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_U67 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n284), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n286), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n285), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n283) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_U66 ( .A(
        Red_StateRegOutput[47]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n270), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n284) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_U65 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n269), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n268), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n267), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n271), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n270) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_U64 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n266), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n276), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n265), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n264), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n263), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n267) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_U63 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n262), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n261), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n280), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n260), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n265) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_U62 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n264), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n276) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_U61 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n275), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n274), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n266) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_U60 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n259), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n268) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_U59 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n258), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n257), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n256), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n269) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_U58 ( .A(
        Red_StateRegOutput[44]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n255), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n285) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_U57 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n254), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n264), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n253), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n252), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n255) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_U56 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n280), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n259), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n251), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n252) );
  NAND4_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_U55 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n256), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n250), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n278), .A4(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n264), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n253) );
  AOI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_U54 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n273), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n249), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n248), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n279), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n254) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_U53 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n260), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n261), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n247), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n279) );
  NOR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_U52 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n280), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n246), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n282), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n248) );
  AND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_U51 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n260), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n261), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n282) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_U50 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n245), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n261) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_U49 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n251), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n271), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n273) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_U48 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n278), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n281), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n259) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_U47 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n264), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n271), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n281) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_U46 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n246), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n258), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n247) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_U45 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n243), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n249), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n258) );
  AND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_U44 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n245), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n244), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n263) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_U43 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n280), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n274), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n244) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_U42 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n251), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n275), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n245) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_U41 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n257), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n275) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_U40 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n251), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n249), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n250) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_U39 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n277), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n257), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n256) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_U38 ( .A(
        Red_StateRegOutput[46]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n242), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n257) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_U37 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n280), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n277) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_U36 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n271), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n246) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_U35 ( .A(
        Red_StateRegOutput[47]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n241), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n271) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_U34 ( .A(
        F_SD2_RedSB_inst_n42), .B(F_SD2_RedSB_inst_n44), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n241) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_U33 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n264), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n243), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n272) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_U32 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n251), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n243) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_U31 ( .A(
        Red_StateRegOutput[45]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n240), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n251) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_U30 ( .A(
        F_SD2_RedSB_inst_n41), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n239), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n264) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_U29 ( .A(
        Red_StateRegOutput[44]), .B(F_SD2_RedSB_inst_n43), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n239) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_U28 ( .A(
        F_SD2_RedSB_inst_n42), .B(F_SD2_RedSB_inst_n43), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n242) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_U27 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n278), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n249), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n260) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_U26 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n274), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n249) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_U25 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n238), .B(
        Red_StateRegOutput[48]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n274) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_U24 ( .A(
        F_SD2_RedSB_inst_n43), .B(F_SD2_RedSB_inst_n44), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n238) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_U23 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n262), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n278) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_U22 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n237), .B(
        Red_StateRegOutput[43]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n262) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_U21 ( .A(
        F_SD2_RedSB_inst_n42), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n240), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n237) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_U20 ( .A(
        F_SD2_RedSB_inst_n41), .B(F_SD2_RedSB_inst_n44), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n240) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_U19 ( .A(
        Red_StateRegOutput[43]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n236), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n289) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_U18 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n260), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n232), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n234), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n235), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n236) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_U17 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n263), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n271), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n263), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n250), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n262), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n235) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_U16 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n245), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n259), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n244), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n259), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n233), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n234) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_U15 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n262), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n247), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n233) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_U14 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n280), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n272), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n246), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n256), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n232) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_U13 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n286), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n288), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n230), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n231), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n289), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n287) );
  OR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_U12 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n285), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n284), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n231) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_U11 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n286), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n230) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_U10 ( .A(
        Red_StateRegOutput[42]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n229), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n280) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_U9 ( .A(
        F_SD2_RedSB_inst_n41), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n242), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n229) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_U8 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n228), .B(
        Red_StateRegOutput[42]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n286) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_U7 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n224), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n279), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n227), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n228) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_U6 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n278), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n225), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n277), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n226), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n227) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_U5 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n276), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n274), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n275), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n226) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_U4 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n271), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n272), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n275), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n273), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n225) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_U3 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n282), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n281), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n280), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_45_n224) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_U73 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n277), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n276), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n279), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n278) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_U72 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n275), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n274), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n273), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n277) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_U71 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n272), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n279) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_U70 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n266), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n265), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n264), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n267) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_U69 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n265), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n269) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_U68 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n280), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n263) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_U67 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n261), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n260), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n280) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_U66 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n264), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n281), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n258), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n276) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_U65 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n283), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n275), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n259) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_U64 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n264), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n257), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n283) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_U63 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n261), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n262), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n254), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n285), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n255) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_U62 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n272), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n253), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n285) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_U61 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n270), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n252), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n282) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_U60 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n286), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n274) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_U59 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n257), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n251), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n286) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_U58 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n250), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n249), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n248), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n256) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_U57 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n260), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n271), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n250), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n248) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_U56 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n273), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n247), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n246), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n249) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_U55 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n284), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n246) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_U54 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n270), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n252), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n284) );
  OR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_U53 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n275), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n253), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n252) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_U52 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n266), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n270) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_U51 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n254), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n275), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n247) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_U50 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n281), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n254) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_U49 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n272), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n244), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n243), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n245) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_U48 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n260), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n262), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n242), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n241), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n243) );
  OR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_U47 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n250), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n271), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n268), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n241) );
  OR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_U46 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n281), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n253), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n261), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n268) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_U45 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n257), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n250) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_U44 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n266), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n251), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n265), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n240), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n253), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n242) );
  AND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_U43 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n266), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n251), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n240) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_U42 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n275), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n257), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n265) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_U41 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n264), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n281), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n251) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_U40 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n261), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n264) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_U39 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n272), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n273), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n266) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_U38 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n273), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n253), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n262) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_U37 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n271), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n273) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_U36 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n275), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n281), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n260) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_U35 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n258), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n275) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_U34 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n258), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n239), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n261), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n239), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n253), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n244) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_U33 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n238), .B(
        Red_StateRegOutput[42]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n253) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_U32 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n237), .B(
        F_SD2_RedSB_inst_n42), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n238) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_U31 ( .A(
        Red_StateRegOutput[44]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n237), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n261) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_U30 ( .A(
        F_SD2_RedSB_inst_n43), .B(F_SD2_RedSB_inst_n41), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n237) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_U29 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n257), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n281), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n271), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n239) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_U28 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n236), .B(
        Red_StateRegOutput[45]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n271) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_U27 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n235), .B(
        F_SD2_RedSB_inst_n42), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n281) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_U26 ( .A(
        Red_StateRegOutput[47]), .B(F_SD2_RedSB_inst_n44), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n235) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_U25 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n234), .B(
        Red_StateRegOutput[43]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n257) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_U24 ( .A(
        F_SD2_RedSB_inst_n42), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n236), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n234) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_U23 ( .A(
        F_SD2_RedSB_inst_n41), .B(F_SD2_RedSB_inst_n44), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n236) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_U22 ( .A(
        Red_StateRegOutput[48]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n233), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n258) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_U21 ( .A(
        F_SD2_RedSB_inst_n43), .B(F_SD2_RedSB_inst_n44), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n233) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_U20 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n232), .B(
        Red_StateRegOutput[46]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n272) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_U19 ( .A(
        F_SD2_RedSB_inst_n43), .B(F_SD2_RedSB_inst_n42), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n232) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_U18 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n217), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n220), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n226), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n230), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n231), .ZN(Red_Feedback[74])
         );
  NOR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_U17 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n220), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n230), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n226), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n231) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_U16 ( .A(
        Red_StateRegOutput[47]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n229), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n230) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_U15 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n285), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n286), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n227), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n228), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n229) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_U14 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n279), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n280), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n278), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n228) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_U13 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n284), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n282), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n284), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n283), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n281), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n227) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_U12 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n224), .B2(
        Red_StateRegOutput[44]), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n225), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n226) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_U11 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n224), .B2(
        Red_StateRegOutput[44]), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n217), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n225) );
  AOI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_U10 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n271), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n221), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n222), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n223), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n224) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_U9 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n262), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n286), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n263), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n271), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n223) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_U8 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n270), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n269), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n267), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n268), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n222) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_U7 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n285), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n259), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n276), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n221) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_U6 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n219), .B(
        Red_StateRegOutput[43]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n220) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_U5 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n218), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n256), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n219) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_U4 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n265), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n255), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n282), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n274), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n218) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_U3 ( .A(
        Red_StateRegOutput[42]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n245), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_46_n217) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_U73 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n284), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n283), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n282), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n281), .ZN(Red_Feedback[75])
         );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_U72 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n280), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n281), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n279), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n283) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_U71 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n280), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n281), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n282), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n279) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_U70 ( .A(
        Red_StateRegOutput[47]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n278), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n282) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_U69 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n277), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n276), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n278) );
  NAND4_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_U68 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n275), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n274), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n273), .A4(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n272), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n276) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_U67 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n271), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n270), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n269), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n268), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n277) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_U66 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n267), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n268) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_U65 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n274), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n266), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n265), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n264), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n270) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_U64 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n263), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n265) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_U63 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n262), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n272), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n261), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n260), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n266) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_U62 ( .A(
        Red_StateRegOutput[43]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n259), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n281) );
  NOR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_U61 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n258), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n257), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n256), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n259) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_U60 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n255), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n254), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n255), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n253), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n252), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n256) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_U59 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n273), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n263), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n252) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_U58 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n251), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n250), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n263) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_U57 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n275), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n262), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n253) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_U56 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n271), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n269), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n254) );
  AOI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_U55 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n275), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n249), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n248), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n247), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n257) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_U54 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n246), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n245), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n275), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n247) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_U53 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n271), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n244), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n249) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_U52 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n245), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n271) );
  NOR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_U51 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n251), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n244), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n250), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n258) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_U50 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n260), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n248), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n250) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_U49 ( .A(
        Red_StateRegOutput[42]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n243), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n280) );
  AOI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_U48 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n275), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n242), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n241), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n240), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n243) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_U47 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n251), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n239), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n255), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n238), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n240) );
  OR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_U46 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n251), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n239), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n260), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n238) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_U45 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n237), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n248), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n244), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n255) );
  NOR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_U44 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n237), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n236), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n272), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n241) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_U43 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n274), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n262), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n246), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n235), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n236) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_U42 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n234), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n260), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n233), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n242) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_U41 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n232), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n246), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n262), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n233) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_U40 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n231), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n234) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_U39 ( .A(
        Red_StateRegOutput[44]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n230), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n284) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_U38 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n262), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n229), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n228), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n230) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_U37 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n267), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n227), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n226), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n264), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n228) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_U36 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n244), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n225), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n264) );
  NAND4_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_U35 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n237), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n269), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n274), .A4(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n227), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n226) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_U34 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n272), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n269) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_U33 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n237), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n273), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n262), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n231), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n267) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_U32 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n245), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n248), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n231) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_U31 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n244), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n239), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n273) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_U30 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n245), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n225), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n239) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_U29 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n260), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n237) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_U28 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n274), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n224), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n223), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n251), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n229) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_U27 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n232), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n244), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n261), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n244), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n235), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n224) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_U26 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n275), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n245), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n235) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_U25 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n227), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n275) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_U24 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n251), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n261) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_U23 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n227), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n272), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n251) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_U22 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n222), .B(
        Red_StateRegOutput[46]), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n272) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_U21 ( .A(
        F_SD2_RedSB_inst_n42), .B(F_SD2_RedSB_inst_n43), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n222) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_U20 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n221), .B(
        Red_StateRegOutput[45]), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n227) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_U19 ( .A(
        F_SD2_RedSB_inst_n41), .B(F_SD2_RedSB_inst_n44), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n221) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_U18 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n246), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n244) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_U17 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n220), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n219), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n246) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_U16 ( .A(
        F_SD2_RedSB_inst_n44), .B(Red_StateRegOutput[43]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n220) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_U15 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n223), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n232) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_U14 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n260), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n245), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n223) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_U13 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n218), .B(
        Red_StateRegOutput[47]), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n245) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_U12 ( .A(
        F_SD2_RedSB_inst_n42), .B(F_SD2_RedSB_inst_n44), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n218) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_U11 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n217), .B(
        F_SD2_RedSB_inst_n43), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n260) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_U10 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n219), .B(
        Red_StateRegOutput[42]), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n217) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_U9 ( .A(
        F_SD2_RedSB_inst_n41), .B(F_SD2_RedSB_inst_n42), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n219) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_U8 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n248), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n274) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_U7 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n216), .B(
        Red_StateRegOutput[48]), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n248) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_U6 ( .A(
        F_SD2_RedSB_inst_n43), .B(F_SD2_RedSB_inst_n44), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n216) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_U5 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n225), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n262) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_U4 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n215), .B(
        F_SD2_RedSB_inst_n43), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n225) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_U3 ( .A(
        Red_StateRegOutput[44]), .B(F_SD2_RedSB_inst_n41), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_47_n215) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_U65 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n283), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n282), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n281), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n280), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n279), .ZN(Red_Feedback[76])
         );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_U64 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n283), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n282), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n281), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n279) );
  MUX2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_U63 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n283), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n282), .S(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n278), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n280) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_U62 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n277), .B(
        Red_StateRegOutput[44]), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n278) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_U61 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n276), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n275), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n274), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n277) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_U60 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n273), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n274) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_U59 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n272), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n271), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n270), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n269), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n268), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n273) );
  AND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_U58 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n267), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n266), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n265), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n269) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_U57 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n266), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n264), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n263), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n262), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n275) );
  AOI222_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_U56 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n261), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n260), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n261), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n259), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n260), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n259), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n263) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_U55 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n258), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n268), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n259) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_U54 ( .A(
        Red_StateRegOutput[42]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n257), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n281) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_U53 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n268), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n256), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n255), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n257) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_U52 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n268), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n254), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n262), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n255) );
  AOI222_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_U51 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n261), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n260), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n261), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n253), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n260), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n253), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n254) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_U50 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n276), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n258), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n253) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_U49 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n252), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n251), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n250), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n249), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n256) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_U48 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n276), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n266), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n248), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n247), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n252) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_U47 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n264), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n247) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_U46 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n272), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n258), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n264) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_U45 ( .A(
        Red_StateRegOutput[43]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n246), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n282) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_U44 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n248), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n262), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n245), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n244), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n246) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_U43 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n248), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n243), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n244) );
  AOI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_U42 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n271), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n242), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n241), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n240), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n245) );
  NOR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_U41 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n270), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n239), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n250), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n240) );
  AND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_U40 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n238), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n268), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n260), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n241) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_U39 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n248), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n266), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n260) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_U38 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n251), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n237), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n249), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n238) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_U37 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n276), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n270), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n249) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_U36 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n258), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n236), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n262) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_U35 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n237), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n258) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_U34 ( .A(
        Red_StateRegOutput[47]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n235), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n283) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_U33 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n234), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n237), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n233), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n237), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n232), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n235) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_U32 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n251), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n268), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n267), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n236), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n271), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n232) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_U31 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n250), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n276), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n271) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_U30 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n237), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n248), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n250) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_U29 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n239), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n272), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n236) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_U28 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n242), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n265), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n243), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n233) );
  AND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_U27 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n261), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n231), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n243) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_U26 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n276), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n248), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n265) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_U25 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n230), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n229), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n248) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_U24 ( .A(
        F_SD2_RedSB_inst_n41), .B(Red_StateRegOutput[43]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n230) );
  OR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_U23 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n261), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n231), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n242) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_U22 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n268), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n266), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n231) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_U21 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n228), .B(
        Red_StateRegOutput[42]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n268) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_U20 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n227), .B(
        F_SD2_RedSB_inst_n42), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n228) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_U19 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n267), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n270), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n261) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_U18 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n272), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n270) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_U17 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n226), .B(
        Red_StateRegOutput[45]), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n272) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_U16 ( .A(
        F_SD2_RedSB_inst_n41), .B(F_SD2_RedSB_inst_n44), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n226) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_U15 ( .A(
        Red_StateRegOutput[47]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n229), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n237) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_U14 ( .A(
        F_SD2_RedSB_inst_n44), .B(F_SD2_RedSB_inst_n42), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n229) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_U13 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n225), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n234) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_U12 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n267), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n239), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n224), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n225) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_U11 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n267), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n239), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n276), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n224) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_U10 ( .A(
        Red_StateRegOutput[44]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n227), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n276) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_U9 ( .A(
        F_SD2_RedSB_inst_n43), .B(F_SD2_RedSB_inst_n41), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n227) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_U8 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n266), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n239) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_U7 ( .A(
        Red_StateRegOutput[48]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n223), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n266) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_U6 ( .A(
        F_SD2_RedSB_inst_n43), .B(F_SD2_RedSB_inst_n44), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n223) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_U5 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n251), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n267) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_U4 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n222), .B(
        Red_StateRegOutput[46]), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n251) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_U3 ( .A(
        F_SD2_RedSB_inst_n43), .B(F_SD2_RedSB_inst_n42), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_48_n222) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_U69 ( .A(
        Red_StateRegOutput[50]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n280), .Z(Red_Feedback[63])
         );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_U68 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n279), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n278), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n280) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_U67 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n277), .B2(
        Red_StateRegOutput[51]), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n276), .C2(
        Red_StateRegOutput[54]), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n275), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n278) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_U66 ( .A1(
        Red_StateRegOutput[51]), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n277), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n276), .B2(
        Red_StateRegOutput[54]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n275) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_U65 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n274), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n273), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n276) );
  AOI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_U64 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n272), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n271), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n270), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n269), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n273) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_U63 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n268), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n267), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n266), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n265), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n264), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n269) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_U62 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n268), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n263), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n262), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n270) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_U61 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n268), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n263), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n261), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n262) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_U60 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n260), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n259), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n258), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n271) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_U59 ( .A(
        Red_StateRegOutput[49]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n257), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n274) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_U58 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n256), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n255), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n254), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n257) );
  OR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_U57 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n267), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n253), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n252), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n254) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_U56 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n251), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n250), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n249), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n252) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_U55 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n250), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n251), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n248), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n253) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_U54 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n247), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n246), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n245), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n244), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n255) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_U53 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n243), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n242), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n241), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n240), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n247) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_U52 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n239), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n238), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n240), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n237), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n236), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n277) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_U51 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n235), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n234), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n233), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n236) );
  AOI222_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_U50 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n251), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n249), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n251), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n232), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n249), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n232), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n234) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_U49 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n242), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n267), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n232) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_U48 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n263), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n246), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n249) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_U47 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n231), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n251) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_U46 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n256), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n230), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n237) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_U45 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n261), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n263), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n229), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n238) );
  NOR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_U44 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n267), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n244), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n259), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n229) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_U43 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n245), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n246), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n259) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_U42 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n268), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n228), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n244) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_U41 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n256), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n267) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_U40 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n242), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n245), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n261) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_U39 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n264), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n260), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n227), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n279) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_U38 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n246), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n226), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n225), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n227) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_U37 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n246), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n224), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n248), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n225) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_U36 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n235), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n248) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_U35 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n242), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n265), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n235) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_U34 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n239), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n228), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n265) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_U33 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n241), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n243), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n256), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n263), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n224) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_U32 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n240), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n245), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n243) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_U31 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n266), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n242), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n241) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_U30 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n272), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n223), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n258), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n226) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_U29 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n231), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n222), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n258) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_U28 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n240), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n228), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n223) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_U27 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n231), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n222), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n260) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_U26 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n228), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n256), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n222) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_U25 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n221), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n220), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n256) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_U24 ( .A(
        Red_StateRegOutput[49]), .B(F_SD2_RedSB_inst_n45), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n221) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_U23 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n263), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n228) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_U22 ( .A(
        Red_StateRegOutput[55]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n219), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n263) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_U21 ( .A(
        F_SD2_RedSB_inst_n48), .B(F_SD2_RedSB_inst_n47), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n219) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_U20 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n239), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n268), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n231) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_U19 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n266), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n268) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_U18 ( .A(
        Red_StateRegOutput[53]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n220), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n266) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_U17 ( .A(
        F_SD2_RedSB_inst_n46), .B(F_SD2_RedSB_inst_n47), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n220) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_U16 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n240), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n239) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_U15 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n218), .B(
        Red_StateRegOutput[52]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n240) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_U14 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n230), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n264) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_U13 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n250), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n246), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n230) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_U12 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n217), .B(
        F_SD2_RedSB_inst_n46), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n246) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_U11 ( .A(
        Red_StateRegOutput[50]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n218), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n217) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_U10 ( .A(
        F_SD2_RedSB_inst_n48), .B(F_SD2_RedSB_inst_n45), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n218) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_U9 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n242), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n245), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n250) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_U8 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n233), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n245) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_U7 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n216), .B(
        Red_StateRegOutput[51]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n233) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_U6 ( .A(
        F_SD2_RedSB_inst_n45), .B(F_SD2_RedSB_inst_n47), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n216) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_U5 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n272), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n242) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_U4 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n215), .B(
        F_SD2_RedSB_inst_n46), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n272) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_U3 ( .A(
        Red_StateRegOutput[54]), .B(F_SD2_RedSB_inst_n48), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_49_n215) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_U67 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n265), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n264), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n270), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n271), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n266) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_U66 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n263), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n262), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n271) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_U65 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n261), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n270), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n260), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n259), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n265) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_U64 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n258), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n270) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_U63 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n272), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n267) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_U62 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n263), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n262), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n272) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_U61 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n274), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n254), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n262) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_U60 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n268), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n255), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n275) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_U59 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n258), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n264), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n255) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_U58 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n269), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n268) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_U57 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n257), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n264), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n253) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_U56 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n277), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n264) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_U55 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n277), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n254), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n251) );
  AND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_U54 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n276), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n273), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n263) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_U53 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n274), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n258), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n260) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_U52 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n256), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n274) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_U51 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n256), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n276), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n261) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_U50 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n257), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n276) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_U49 ( .A(
        Red_StateRegOutput[54]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n250), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n277) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_U48 ( .A(
        F_SD2_RedSB_inst_n47), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n249), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n269) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_U47 ( .A(
        Red_StateRegOutput[51]), .B(F_SD2_RedSB_inst_n45), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n249) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_U46 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n273), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n252), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n259) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_U45 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n254), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n252) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_U44 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n248), .B(
        Red_StateRegOutput[49]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n254) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_U43 ( .A(
        F_SD2_RedSB_inst_n45), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n247), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n248) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_U42 ( .A(
        Red_StateRegOutput[53]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n247), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n273) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_U41 ( .A(
        F_SD2_RedSB_inst_n47), .B(F_SD2_RedSB_inst_n46), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n247) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_U40 ( .A(
        Red_StateRegOutput[55]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n246), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n256) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_U39 ( .A(
        F_SD2_RedSB_inst_n47), .B(F_SD2_RedSB_inst_n48), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n246) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_U38 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n245), .B(
        Red_StateRegOutput[52]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n257) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_U37 ( .A(
        F_SD2_RedSB_inst_n45), .B(F_SD2_RedSB_inst_n48), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n245) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_U36 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n244), .B(
        Red_StateRegOutput[50]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n258) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_U35 ( .A(
        F_SD2_RedSB_inst_n45), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n250), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n244) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_U34 ( .A(
        F_SD2_RedSB_inst_n46), .B(F_SD2_RedSB_inst_n48), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n250) );
  AOI222_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_U33 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n221), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n230), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n221), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n238), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n230), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n243), .ZN(Red_Feedback[64])
         );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_U32 ( .A(
        Red_StateRegOutput[50]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n242), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n243) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_U31 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n255), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n239), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n240), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n241), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n242) );
  NAND4_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_U30 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n254), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n257), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n268), .A4(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n260), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n241) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_U29 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n275), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n267), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n266), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n240) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_U28 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n226), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n239) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_U27 ( .A(
        Red_StateRegOutput[54]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n237), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n238) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_U26 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n277), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n234), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n275), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n236), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n237) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_U25 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n276), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n232), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n235), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n236) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_U24 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n259), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n235) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_U23 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n272), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n231), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n271), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n233), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n234) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_U22 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n273), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n274), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n268), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n232), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n233) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_U21 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n273), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n274), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n232) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_U20 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n270), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n269), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n231) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_U19 ( .A(
        Red_StateRegOutput[51]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n229), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n230) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_U18 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n252), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n222), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n225), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n228), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n229) );
  NAND4_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_U17 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n269), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n259), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n226), .A4(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n227), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n228) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_U16 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n258), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n227) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_U15 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n256), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n257), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n226) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_U14 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n224), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n260), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n224), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n251), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n268), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n225) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_U13 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n215), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n223), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n224) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_U12 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n256), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n253), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n263), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n251), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n223) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_U11 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n257), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n275), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n222) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_U10 ( .A(
        Red_StateRegOutput[49]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n220), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n221) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_U9 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n254), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n218), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n219), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n220) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_U8 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n254), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n215), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n214), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n219) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_U7 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n255), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n216), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n273), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n217), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n218) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_U6 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n258), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n253), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n268), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n274), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n217) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_U5 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n257), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n268), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n216) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_U4 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n277), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n261), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n263), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n260), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n215) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_U3 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n263), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n260), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n264), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n269), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_50_n214) );
  MUX2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_U54 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n240), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n239), .S(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n238), .Z(Red_Feedback[65])
         );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_U53 ( .A(
        Red_StateRegOutput[51]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n237), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n238) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_U52 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n236), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n235), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n234), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n233), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n237) );
  OR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_U51 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n232), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n231), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n230), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n233) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_U50 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n229), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n228), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n227), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n234) );
  AOI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_U49 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n226), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n225), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n224), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n223), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n236) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_U48 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n222), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n221), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n220), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n221), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n219), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n223) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_U47 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n226), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n225), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n218), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n221) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_U46 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n217), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n216), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n225) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_U45 ( .A(
        Red_StateRegOutput[54]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n215), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n239) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_U44 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n214), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n230), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n213), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n212), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n215) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_U43 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n228), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n226), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n211), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n232), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n212) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_U42 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n210), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n228), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n210), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n226), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n216), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n213) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_U41 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n220), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n216) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_U40 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n209), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n226) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_U39 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n208), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n207), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n228) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_U38 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n219), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n206), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n205), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n210) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_U37 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n219), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n206), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n208), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n205) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_U36 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n235), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n208) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_U35 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n222), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n204), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n229), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n214) );
  AND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_U34 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n206), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n219), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n204) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_U33 ( .A(
        Red_StateRegOutput[50]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n203), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n240) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_U32 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n202), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n201), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n200), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n201), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n199), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n203) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_U31 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n198), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n197), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n230), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n209), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n199) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_U30 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n227), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n220), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n218), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n197) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_U29 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n207), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n218) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_U28 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n222), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n201), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n227) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_U27 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n198), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n230), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n209), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n230), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n217), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n200) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_U26 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n231), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n206), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n209) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_U25 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n207), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n235), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n220), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n230) );
  AOI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_U24 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n229), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n211), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n207), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n224), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n198) );
  NOR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_U23 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n231), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n220), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n201), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n224) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_U22 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n219), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n220), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n211) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_U21 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n196), .B(
        Red_StateRegOutput[54]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n220) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_U20 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n201), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n219) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_U19 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n232), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n206), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n229) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_U18 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n195), .B(
        Red_StateRegOutput[53]), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n206) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_U17 ( .A(
        F_SD2_RedSB_inst_n47), .B(F_SD2_RedSB_inst_n46), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n195) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_U16 ( .A(
        Red_StateRegOutput[55]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n194), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n201) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_U15 ( .A(
        F_SD2_RedSB_inst_n47), .B(F_SD2_RedSB_inst_n48), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n194) );
  NOR4_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_U14 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n207), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n231), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n232), .A4(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n235), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n202) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_U13 ( .A(
        Red_StateRegOutput[51]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n193), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n235) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_U12 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n217), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n232) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_U11 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n192), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n193), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n217) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_U10 ( .A(
        F_SD2_RedSB_inst_n45), .B(F_SD2_RedSB_inst_n47), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n193) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_U9 ( .A(
        F_SD2_RedSB_inst_n46), .B(Red_StateRegOutput[49]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n192) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_U8 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n222), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n231) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_U7 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n191), .B(
        Red_StateRegOutput[52]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n222) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_U6 ( .A(
        F_SD2_RedSB_inst_n45), .B(F_SD2_RedSB_inst_n48), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n191) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_U5 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n190), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n196), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n207) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_U4 ( .A(
        F_SD2_RedSB_inst_n46), .B(F_SD2_RedSB_inst_n48), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n196) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_U3 ( .A(
        F_SD2_RedSB_inst_n45), .B(Red_StateRegOutput[50]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_51_n190) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_U71 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n288), .B(
        Red_StateRegOutput[49]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n291) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_U70 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n287), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n286), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n288) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_U69 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n285), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n284), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n283), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n282), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n286) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_U68 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n281), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n282) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_U67 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n280), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n279), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n278), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n277), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n287) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_U66 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n276), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n275), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n274), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n277) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_U65 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n273), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n275), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n272), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n271), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n280) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_U64 ( .A(
        Red_StateRegOutput[54]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n270), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n289) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_U63 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n269), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n268), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n267), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n271), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n270) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_U62 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n266), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n276), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n265), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n264), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n263), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n267) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_U61 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n262), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n261), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n283), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n260), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n265) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_U60 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n264), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n276) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_U59 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n275), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n274), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n266) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_U58 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n259), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n268) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_U57 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n258), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n257), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n256), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n269) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_U56 ( .A(
        Red_StateRegOutput[51]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n255), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n290) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_U55 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n254), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n264), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n253), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n252), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n255) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_U54 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n283), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n259), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n251), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n252) );
  NAND4_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_U53 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n256), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n250), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n279), .A4(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n264), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n253) );
  AOI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_U52 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n273), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n249), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n248), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n281), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n254) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_U51 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n260), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n261), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n247), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n281) );
  NOR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_U50 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n283), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n246), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n285), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n248) );
  AND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_U49 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n260), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n261), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n285) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_U48 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n245), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n261) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_U47 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n251), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n271), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n273) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_U46 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n245), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n243), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n259), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n244) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_U45 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n279), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n284), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n259) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_U44 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n264), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n271), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n284) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_U43 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n246), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n258), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n247) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_U42 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n242), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n249), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n258) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_U41 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n271), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n250), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n263), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n241) );
  AND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_U40 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n245), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n243), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n263) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_U39 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n283), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n274), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n243) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_U38 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n251), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n275), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n245) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_U37 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n257), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n275) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_U36 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n251), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n249), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n250) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_U35 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n278), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n257), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n256) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_U34 ( .A(
        Red_StateRegOutput[53]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n240), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n257) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_U33 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n283), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n278) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_U32 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n271), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n246) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_U31 ( .A(
        Red_StateRegOutput[54]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n239), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n271) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_U30 ( .A(
        F_SD2_RedSB_inst_n46), .B(F_SD2_RedSB_inst_n48), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n239) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_U29 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n264), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n242), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n272) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_U28 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n251), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n242) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_U27 ( .A(
        Red_StateRegOutput[52]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n238), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n251) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_U26 ( .A(
        F_SD2_RedSB_inst_n45), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n237), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n264) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_U25 ( .A(
        Red_StateRegOutput[51]), .B(F_SD2_RedSB_inst_n47), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n237) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_U24 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n236), .B(
        F_SD2_RedSB_inst_n45), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n283) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_U23 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n235), .B(
        Red_StateRegOutput[49]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n236) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_U22 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n240), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n235) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_U21 ( .A(
        F_SD2_RedSB_inst_n46), .B(F_SD2_RedSB_inst_n47), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n240) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_U20 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n279), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n249), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n260) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_U19 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n274), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n249) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_U18 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n234), .B(
        Red_StateRegOutput[55]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n274) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_U17 ( .A(
        F_SD2_RedSB_inst_n47), .B(F_SD2_RedSB_inst_n48), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n234) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_U16 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n262), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n279) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_U15 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n233), .B(
        Red_StateRegOutput[50]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n262) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_U14 ( .A(
        F_SD2_RedSB_inst_n46), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n238), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n233) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_U13 ( .A(
        F_SD2_RedSB_inst_n45), .B(F_SD2_RedSB_inst_n48), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n238) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_U12 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n230), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n228), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n231), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n232), .ZN(Red_Feedback[66])
         );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_U11 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n230), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n224), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n228), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n232) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_U10 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n290), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n289), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n291), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n231) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_U9 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n290), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n289), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n229), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n230) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_U8 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n289), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n291), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n290), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n229) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_U7 ( .A(
        Red_StateRegOutput[50]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n227), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n228) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_U6 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n260), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n225), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n244), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n226), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n227) );
  MUX2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_U5 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n247), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n241), .S(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n262), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n226) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_U4 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n246), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n256), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n272), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n283), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n225) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_U3 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n291), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_52_n224) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_U74 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n287), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n286), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n285), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n284), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n283), .ZN(Red_Feedback[67])
         );
  NOR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_U73 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n286), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n284), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n285), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n283) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_U72 ( .A(
        Red_StateRegOutput[54]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n282), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n284) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_U71 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n281), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n280), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n279), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n278), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n282) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_U70 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n277), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n276), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n277), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n275), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n274), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n278) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_U69 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n273), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n272), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n271), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n279) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_U68 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n270), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n269), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n272), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n271) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_U67 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n268), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n267), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n266), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n270) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_U66 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n265), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n272) );
  AOI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_U65 ( .C1(
        Red_StateRegOutput[51]), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n264), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n263), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n262), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n285) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_U64 ( .A1(
        Red_StateRegOutput[51]), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n264), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n262) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_U63 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n287), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n263) );
  AOI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_U62 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n261), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n260), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n259), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n258), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n264) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_U61 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n257), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n256), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n255), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n254), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n258) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_U60 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n253), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n252), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n251), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n254) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_U59 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n252), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n256) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_U58 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n250), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n261), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n281), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n249), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n259) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_U57 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n273), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n250) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_U56 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n248), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n247), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n273) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_U55 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n280), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n246), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n269), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n260) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_U54 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n251), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n274), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n245), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n269) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_U53 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n276), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n268), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n246) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_U52 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n251), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n244), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n276) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_U51 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n243), .B(
        Red_StateRegOutput[50]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n286) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_U50 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n242), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n241), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n243) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_U49 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n267), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n275), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n252), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n240), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n241) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_U48 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n248), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n249), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n239), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n280), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n240) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_U47 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n265), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n238), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n280) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_U46 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n257), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n237), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n275) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_U45 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n281), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n267) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_U44 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n244), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n236), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n281) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_U43 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n235), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n234), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n233), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n242) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_U42 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n247), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n261), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n235), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n233) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_U41 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n266), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n232), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n231), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n234) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_U40 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n277), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n231) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_U39 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n257), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n237), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n277) );
  OR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_U38 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n268), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n238), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n237) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_U37 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n253), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n257) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_U36 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n239), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n268), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n232) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_U35 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n274), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n239) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_U34 ( .A(
        Red_StateRegOutput[49]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n230), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n287) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_U33 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n265), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n229), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n228), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n230) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_U32 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n247), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n249), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n227), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n226), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n228) );
  OR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_U31 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n235), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n261), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n255), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n226) );
  OR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_U30 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n274), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n238), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n248), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n255) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_U29 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n244), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n235) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_U28 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n253), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n236), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n252), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n225), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n238), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n227) );
  AND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_U27 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n253), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n236), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n225) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_U26 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n268), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n244), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n252) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_U25 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n251), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n274), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n236) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_U24 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n248), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n251) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_U23 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n265), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n266), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n253) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_U22 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n266), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n238), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n249) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_U21 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n261), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n266) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_U20 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n268), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n274), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n247) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_U19 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n245), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n268) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_U18 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n245), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n224), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n248), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n224), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n238), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n229) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_U17 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n223), .B(
        Red_StateRegOutput[49]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n238) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_U16 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n222), .B(
        F_SD2_RedSB_inst_n46), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n223) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_U15 ( .A(
        Red_StateRegOutput[51]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n222), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n248) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_U14 ( .A(
        F_SD2_RedSB_inst_n47), .B(F_SD2_RedSB_inst_n45), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n222) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_U13 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n244), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n274), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n261), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n224) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_U12 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n221), .B(
        Red_StateRegOutput[52]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n261) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_U11 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n220), .B(
        F_SD2_RedSB_inst_n46), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n274) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_U10 ( .A(
        Red_StateRegOutput[54]), .B(F_SD2_RedSB_inst_n48), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n220) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_U9 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n219), .B(
        Red_StateRegOutput[50]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n244) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_U8 ( .A(
        F_SD2_RedSB_inst_n46), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n221), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n219) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_U7 ( .A(
        F_SD2_RedSB_inst_n45), .B(F_SD2_RedSB_inst_n48), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n221) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_U6 ( .A(
        Red_StateRegOutput[55]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n218), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n245) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_U5 ( .A(
        F_SD2_RedSB_inst_n47), .B(F_SD2_RedSB_inst_n48), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n218) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_U4 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n217), .B(
        Red_StateRegOutput[53]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n265) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_U3 ( .A(
        F_SD2_RedSB_inst_n47), .B(F_SD2_RedSB_inst_n46), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_53_n217) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_U73 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n284), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n283), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n282), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n281), .ZN(Red_Feedback[68])
         );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_U72 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n280), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n281), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n279), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n283) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_U71 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n280), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n281), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n282), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n279) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_U70 ( .A(
        Red_StateRegOutput[54]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n278), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n282) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_U69 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n277), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n276), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n278) );
  NAND4_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_U68 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n275), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n274), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n273), .A4(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n272), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n276) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_U67 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n271), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n270), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n269), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n268), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n277) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_U66 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n267), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n268) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_U65 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n274), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n266), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n265), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n264), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n270) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_U64 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n263), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n265) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_U63 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n262), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n272), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n261), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n260), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n266) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_U62 ( .A(
        Red_StateRegOutput[50]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n259), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n281) );
  NOR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_U61 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n258), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n257), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n256), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n259) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_U60 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n255), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n254), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n255), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n253), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n252), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n256) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_U59 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n273), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n263), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n252) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_U58 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n251), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n250), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n263) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_U57 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n275), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n262), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n253) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_U56 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n271), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n269), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n254) );
  AOI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_U55 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n275), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n249), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n248), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n247), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n257) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_U54 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n246), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n245), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n275), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n247) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_U53 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n271), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n244), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n249) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_U52 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n245), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n271) );
  NOR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_U51 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n251), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n244), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n250), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n258) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_U50 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n260), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n248), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n250) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_U49 ( .A(
        Red_StateRegOutput[49]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n243), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n280) );
  AOI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_U48 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n275), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n242), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n241), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n240), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n243) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_U47 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n251), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n239), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n255), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n238), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n240) );
  OR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_U46 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n251), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n239), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n260), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n238) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_U45 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n237), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n248), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n244), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n255) );
  NOR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_U44 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n237), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n236), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n272), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n241) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_U43 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n274), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n262), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n246), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n235), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n236) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_U42 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n234), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n260), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n233), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n242) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_U41 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n232), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n246), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n262), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n233) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_U40 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n231), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n234) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_U39 ( .A(
        Red_StateRegOutput[51]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n230), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n284) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_U38 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n262), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n229), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n228), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n230) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_U37 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n267), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n227), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n226), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n264), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n228) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_U36 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n244), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n225), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n264) );
  NAND4_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_U35 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n237), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n269), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n274), .A4(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n227), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n226) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_U34 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n272), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n269) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_U33 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n237), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n273), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n262), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n231), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n267) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_U32 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n245), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n248), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n231) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_U31 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n244), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n239), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n273) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_U30 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n245), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n225), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n239) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_U29 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n260), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n237) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_U28 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n274), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n224), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n223), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n251), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n229) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_U27 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n232), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n244), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n261), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n244), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n235), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n224) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_U26 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n275), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n245), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n235) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_U25 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n227), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n275) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_U24 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n251), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n261) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_U23 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n227), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n272), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n251) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_U22 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n222), .B(
        Red_StateRegOutput[53]), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n272) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_U21 ( .A(
        F_SD2_RedSB_inst_n46), .B(F_SD2_RedSB_inst_n47), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n222) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_U20 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n221), .B(
        Red_StateRegOutput[52]), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n227) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_U19 ( .A(
        F_SD2_RedSB_inst_n45), .B(F_SD2_RedSB_inst_n48), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n221) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_U18 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n246), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n244) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_U17 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n220), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n219), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n246) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_U16 ( .A(
        F_SD2_RedSB_inst_n48), .B(Red_StateRegOutput[50]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n220) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_U15 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n223), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n232) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_U14 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n260), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n245), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n223) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_U13 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n218), .B(
        Red_StateRegOutput[54]), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n245) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_U12 ( .A(
        F_SD2_RedSB_inst_n46), .B(F_SD2_RedSB_inst_n48), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n218) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_U11 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n217), .B(
        F_SD2_RedSB_inst_n47), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n260) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_U10 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n219), .B(
        Red_StateRegOutput[49]), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n217) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_U9 ( .A(
        F_SD2_RedSB_inst_n45), .B(F_SD2_RedSB_inst_n46), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n219) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_U8 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n248), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n274) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_U7 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n216), .B(
        Red_StateRegOutput[55]), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n248) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_U6 ( .A(
        F_SD2_RedSB_inst_n47), .B(F_SD2_RedSB_inst_n48), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n216) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_U5 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n225), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n262) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_U4 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n215), .B(
        F_SD2_RedSB_inst_n47), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n225) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_U3 ( .A(
        Red_StateRegOutput[51]), .B(F_SD2_RedSB_inst_n45), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_54_n215) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_U65 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n283), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n282), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n281), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n280), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n279), .ZN(Red_Feedback[69])
         );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_U64 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n283), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n282), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n281), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n279) );
  MUX2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_U63 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n283), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n282), .S(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n278), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n280) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_U62 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n277), .B(
        Red_StateRegOutput[51]), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n278) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_U61 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n276), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n275), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n274), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n277) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_U60 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n273), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n274) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_U59 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n272), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n271), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n270), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n269), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n268), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n273) );
  AND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_U58 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n267), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n266), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n265), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n269) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_U57 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n266), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n264), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n263), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n262), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n275) );
  AOI222_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_U56 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n261), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n260), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n261), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n259), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n260), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n259), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n263) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_U55 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n258), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n268), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n259) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_U54 ( .A(
        Red_StateRegOutput[49]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n257), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n281) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_U53 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n268), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n256), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n255), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n257) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_U52 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n268), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n254), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n262), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n255) );
  AOI222_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_U51 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n261), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n260), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n261), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n253), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n260), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n253), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n254) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_U50 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n276), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n258), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n253) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_U49 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n252), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n251), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n250), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n249), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n256) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_U48 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n276), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n266), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n248), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n247), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n252) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_U47 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n264), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n247) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_U46 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n272), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n258), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n264) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_U45 ( .A(
        Red_StateRegOutput[50]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n246), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n282) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_U44 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n248), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n262), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n245), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n244), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n246) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_U43 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n248), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n243), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n244) );
  AOI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_U42 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n271), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n242), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n241), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n240), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n245) );
  NOR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_U41 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n270), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n239), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n250), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n240) );
  AND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_U40 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n238), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n268), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n260), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n241) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_U39 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n248), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n266), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n260) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_U38 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n251), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n237), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n249), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n238) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_U37 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n276), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n270), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n249) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_U36 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n258), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n236), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n262) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_U35 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n237), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n258) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_U34 ( .A(
        Red_StateRegOutput[54]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n235), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n283) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_U33 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n234), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n237), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n233), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n237), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n232), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n235) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_U32 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n251), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n268), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n267), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n236), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n271), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n232) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_U31 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n250), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n276), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n271) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_U30 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n237), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n248), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n250) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_U29 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n239), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n272), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n236) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_U28 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n242), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n265), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n243), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n233) );
  AND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_U27 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n261), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n231), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n243) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_U26 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n276), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n248), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n265) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_U25 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n230), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n229), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n248) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_U24 ( .A(
        F_SD2_RedSB_inst_n45), .B(Red_StateRegOutput[50]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n230) );
  OR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_U23 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n261), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n231), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n242) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_U22 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n268), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n266), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n231) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_U21 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n228), .B(
        Red_StateRegOutput[49]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n268) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_U20 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n227), .B(
        F_SD2_RedSB_inst_n46), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n228) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_U19 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n267), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n270), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n261) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_U18 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n272), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n270) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_U17 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n226), .B(
        Red_StateRegOutput[52]), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n272) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_U16 ( .A(
        F_SD2_RedSB_inst_n45), .B(F_SD2_RedSB_inst_n48), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n226) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_U15 ( .A(
        Red_StateRegOutput[54]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n229), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n237) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_U14 ( .A(
        F_SD2_RedSB_inst_n48), .B(F_SD2_RedSB_inst_n46), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n229) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_U13 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n225), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n234) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_U12 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n267), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n239), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n224), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n225) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_U11 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n267), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n239), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n276), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n224) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_U10 ( .A(
        Red_StateRegOutput[51]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n227), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n276) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_U9 ( .A(
        F_SD2_RedSB_inst_n47), .B(F_SD2_RedSB_inst_n45), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n227) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_U8 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n266), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n239) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_U7 ( .A(
        Red_StateRegOutput[55]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n223), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n266) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_U6 ( .A(
        F_SD2_RedSB_inst_n47), .B(F_SD2_RedSB_inst_n48), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n223) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_U5 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n251), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n267) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_U4 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n222), .B(
        Red_StateRegOutput[53]), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n251) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_U3 ( .A(
        F_SD2_RedSB_inst_n47), .B(F_SD2_RedSB_inst_n46), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_55_n222) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_U69 ( .A(
        Red_StateRegOutput[57]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n280), .Z(Red_Feedback[28])
         );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_U68 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n279), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n278), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n280) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_U67 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n277), .B2(
        Red_StateRegOutput[58]), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n276), .C2(
        Red_StateRegOutput[61]), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n275), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n278) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_U66 ( .A1(
        Red_StateRegOutput[58]), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n277), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n276), .B2(
        Red_StateRegOutput[61]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n275) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_U65 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n274), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n273), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n276) );
  AOI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_U64 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n272), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n271), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n270), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n269), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n273) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_U63 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n268), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n267), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n266), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n265), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n264), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n269) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_U62 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n268), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n263), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n262), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n270) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_U61 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n268), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n263), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n261), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n262) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_U60 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n260), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n259), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n258), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n271) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_U59 ( .A(
        Red_StateRegOutput[56]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n257), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n274) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_U58 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n256), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n255), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n254), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n257) );
  OR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_U57 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n267), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n253), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n252), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n254) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_U56 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n251), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n250), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n249), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n252) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_U55 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n250), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n251), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n248), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n253) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_U54 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n247), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n246), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n245), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n244), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n255) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_U53 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n243), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n242), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n241), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n240), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n247) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_U52 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n239), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n238), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n240), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n237), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n236), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n277) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_U51 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n235), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n234), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n233), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n236) );
  AOI222_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_U50 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n251), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n249), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n251), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n232), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n249), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n232), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n234) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_U49 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n242), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n267), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n232) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_U48 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n263), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n246), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n249) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_U47 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n231), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n251) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_U46 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n256), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n230), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n237) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_U45 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n261), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n263), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n229), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n238) );
  NOR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_U44 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n267), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n244), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n259), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n229) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_U43 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n245), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n246), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n259) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_U42 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n268), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n228), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n244) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_U41 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n256), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n267) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_U40 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n242), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n245), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n261) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_U39 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n264), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n260), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n227), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n279) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_U38 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n246), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n226), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n225), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n227) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_U37 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n246), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n224), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n248), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n225) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_U36 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n235), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n248) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_U35 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n242), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n265), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n235) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_U34 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n239), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n228), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n265) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_U33 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n241), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n243), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n256), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n263), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n224) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_U32 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n240), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n245), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n243) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_U31 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n266), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n242), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n241) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_U30 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n272), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n223), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n258), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n226) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_U29 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n231), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n222), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n258) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_U28 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n240), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n228), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n223) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_U27 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n231), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n222), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n260) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_U26 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n228), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n256), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n222) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_U25 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n221), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n220), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n256) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_U24 ( .A(
        Red_StateRegOutput[56]), .B(F_SD2_RedSB_inst_n49), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n221) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_U23 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n263), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n228) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_U22 ( .A(
        Red_StateRegOutput[62]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n219), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n263) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_U21 ( .A(
        F_SD2_RedSB_inst_n52), .B(F_SD2_RedSB_inst_n51), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n219) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_U20 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n239), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n268), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n231) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_U19 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n266), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n268) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_U18 ( .A(
        Red_StateRegOutput[60]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n220), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n266) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_U17 ( .A(
        F_SD2_RedSB_inst_n50), .B(F_SD2_RedSB_inst_n51), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n220) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_U16 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n240), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n239) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_U15 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n218), .B(
        Red_StateRegOutput[59]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n240) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_U14 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n230), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n264) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_U13 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n250), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n246), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n230) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_U12 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n217), .B(
        F_SD2_RedSB_inst_n50), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n246) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_U11 ( .A(
        Red_StateRegOutput[57]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n218), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n217) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_U10 ( .A(
        F_SD2_RedSB_inst_n52), .B(F_SD2_RedSB_inst_n49), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n218) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_U9 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n242), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n245), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n250) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_U8 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n233), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n245) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_U7 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n216), .B(
        Red_StateRegOutput[58]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n233) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_U6 ( .A(
        F_SD2_RedSB_inst_n49), .B(F_SD2_RedSB_inst_n51), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n216) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_U5 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n272), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n242) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_U4 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n215), .B(
        F_SD2_RedSB_inst_n50), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n272) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_U3 ( .A(
        Red_StateRegOutput[61]), .B(F_SD2_RedSB_inst_n52), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_56_n215) );
  AOI222_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_U69 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n279), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n278), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n279), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n277), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n278), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n276), .ZN(Red_Feedback[29])
         );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_U68 ( .A(
        Red_StateRegOutput[61]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n275), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n276) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_U67 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n274), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n273), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n272), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n273), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n271), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n275) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_U66 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n270), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n269), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n268), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n269), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n267), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n271) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_U65 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n266), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n267) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_U64 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n265), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n264), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n268) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_U63 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n263), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n262), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n261), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n272) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_U62 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n260), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n259), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n262) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_U61 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n265), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n264), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n258), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n274) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_U60 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n265), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n264), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n257), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n258) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_U59 ( .A(
        Red_StateRegOutput[57]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n256), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n277) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_U58 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n255), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n254), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n253), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n256) );
  AOI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_U57 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n266), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n252), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n251), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n250), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n253) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_U56 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n249), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n248), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n260), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n261), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n250) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_U55 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n247), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n246), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n261) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_U54 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n245), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n260), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n244), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n243), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n249) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_U53 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n242), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n260) );
  NOR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_U52 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n241), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n240), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n239), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n251) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_U51 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n263), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n252) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_U50 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n247), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n246), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n263) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_U49 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n265), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n238), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n246) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_U48 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n244), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n238), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n254) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_U47 ( .A(
        Red_StateRegOutput[56]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n237), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n278) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_U46 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n238), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n236), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n235), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n237) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_U45 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n238), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n234), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n233), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n235) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_U44 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n244), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n247), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n259), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n248), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n233) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_U43 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n232), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n264), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n239), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n255), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n236) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_U42 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n257), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n241), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n255) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_U41 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n257), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n265), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n242), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n231), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n232) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_U40 ( .A(
        Red_StateRegOutput[58]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n230), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n279) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_U39 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n229), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n259), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n228), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n257), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n227), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n230) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_U38 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n226), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n225), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n224), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n223), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n227) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_U37 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n257), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n244), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n223) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_U36 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n222), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n224) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_U35 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n241), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n266), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n225) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_U34 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n257), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n239), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n266) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_U33 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n242), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n248), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n239) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_U32 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n259), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n257) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_U31 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n234), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n221), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n228) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_U30 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n222), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n247), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n231), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n240), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n221) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_U29 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n241), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n248), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n231) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_U28 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n273), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n248) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_U27 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n273), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n238), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n222) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_U26 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n273), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n245), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n244), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n247), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n234) );
  AND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_U25 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n270), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n264), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n247) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_U24 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n265), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n242), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n244) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_U23 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n240), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n265) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_U22 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n240), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n270), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n245) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_U21 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n241), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n270) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_U20 ( .A(
        Red_StateRegOutput[61]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n220), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n273) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_U19 ( .A(
        F_SD2_RedSB_inst_n51), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n219), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n259) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_U18 ( .A(
        Red_StateRegOutput[58]), .B(F_SD2_RedSB_inst_n49), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n219) );
  NOR4_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_U17 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n242), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n241), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n240), .A4(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n269), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n229) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_U16 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n243), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n269) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_U15 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n264), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n226), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n243) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_U14 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n238), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n226) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_U13 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n218), .B(
        Red_StateRegOutput[56]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n238) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_U12 ( .A(
        F_SD2_RedSB_inst_n49), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n217), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n218) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_U11 ( .A(
        Red_StateRegOutput[60]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n217), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n264) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_U10 ( .A(
        F_SD2_RedSB_inst_n51), .B(F_SD2_RedSB_inst_n50), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n217) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_U9 ( .A(
        Red_StateRegOutput[62]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n216), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n240) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_U8 ( .A(
        F_SD2_RedSB_inst_n51), .B(F_SD2_RedSB_inst_n52), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n216) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_U7 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n215), .B(
        Red_StateRegOutput[59]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n241) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_U6 ( .A(
        F_SD2_RedSB_inst_n49), .B(F_SD2_RedSB_inst_n52), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n215) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_U5 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n214), .B(
        Red_StateRegOutput[57]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n242) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_U4 ( .A(
        F_SD2_RedSB_inst_n49), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n220), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n214) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_U3 ( .A(
        F_SD2_RedSB_inst_n50), .B(F_SD2_RedSB_inst_n52), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_57_n220) );
  MUX2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_U54 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n240), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n239), .S(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n238), .Z(Red_Feedback[30])
         );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_U53 ( .A(
        Red_StateRegOutput[58]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n237), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n238) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_U52 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n236), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n235), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n234), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n233), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n237) );
  OR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_U51 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n232), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n231), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n230), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n233) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_U50 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n229), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n228), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n227), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n234) );
  AOI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_U49 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n226), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n225), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n224), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n223), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n236) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_U48 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n222), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n221), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n220), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n221), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n219), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n223) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_U47 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n226), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n225), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n218), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n221) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_U46 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n217), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n216), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n225) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_U45 ( .A(
        Red_StateRegOutput[61]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n215), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n239) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_U44 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n214), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n230), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n213), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n212), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n215) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_U43 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n228), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n226), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n211), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n232), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n212) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_U42 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n210), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n228), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n210), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n226), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n216), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n213) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_U41 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n220), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n216) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_U40 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n209), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n226) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_U39 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n208), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n207), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n228) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_U38 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n219), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n206), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n205), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n210) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_U37 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n219), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n206), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n208), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n205) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_U36 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n235), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n208) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_U35 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n222), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n204), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n229), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n214) );
  AND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_U34 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n206), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n219), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n204) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_U33 ( .A(
        Red_StateRegOutput[57]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n203), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n240) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_U32 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n202), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n201), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n200), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n201), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n199), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n203) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_U31 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n198), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n197), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n230), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n209), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n199) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_U30 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n227), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n220), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n218), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n197) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_U29 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n207), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n218) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_U28 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n222), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n201), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n227) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_U27 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n198), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n230), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n209), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n230), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n217), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n200) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_U26 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n231), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n206), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n209) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_U25 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n207), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n235), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n220), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n230) );
  AOI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_U24 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n229), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n211), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n207), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n224), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n198) );
  NOR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_U23 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n231), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n220), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n201), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n224) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_U22 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n219), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n220), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n211) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_U21 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n196), .B(
        Red_StateRegOutput[61]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n220) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_U20 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n201), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n219) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_U19 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n232), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n206), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n229) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_U18 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n195), .B(
        Red_StateRegOutput[60]), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n206) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_U17 ( .A(
        F_SD2_RedSB_inst_n51), .B(F_SD2_RedSB_inst_n50), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n195) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_U16 ( .A(
        Red_StateRegOutput[62]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n194), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n201) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_U15 ( .A(
        F_SD2_RedSB_inst_n51), .B(F_SD2_RedSB_inst_n52), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n194) );
  NOR4_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_U14 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n207), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n231), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n232), .A4(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n235), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n202) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_U13 ( .A(
        Red_StateRegOutput[58]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n193), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n235) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_U12 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n217), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n232) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_U11 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n192), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n193), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n217) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_U10 ( .A(
        F_SD2_RedSB_inst_n49), .B(F_SD2_RedSB_inst_n51), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n193) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_U9 ( .A(
        F_SD2_RedSB_inst_n50), .B(Red_StateRegOutput[56]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n192) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_U8 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n222), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n231) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_U7 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n191), .B(
        Red_StateRegOutput[59]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n222) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_U6 ( .A(
        F_SD2_RedSB_inst_n49), .B(F_SD2_RedSB_inst_n52), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n191) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_U5 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n190), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n196), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n207) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_U4 ( .A(
        F_SD2_RedSB_inst_n50), .B(F_SD2_RedSB_inst_n52), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n196) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_U3 ( .A(
        F_SD2_RedSB_inst_n49), .B(Red_StateRegOutput[57]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_58_n190) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_U71 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n289), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n291), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n290), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n288) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_U70 ( .A(
        Red_StateRegOutput[61]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n275), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n289) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_U69 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n274), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n273), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n272), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n276), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n275) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_U68 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n271), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n281), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n270), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n269), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n268), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n272) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_U67 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n267), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n266), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n285), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n265), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n270) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_U66 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n269), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n281) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_U65 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n280), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n279), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n271) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_U64 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n264), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n273) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_U63 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n263), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n262), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n261), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n274) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_U62 ( .A(
        Red_StateRegOutput[58]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n260), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n290) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_U61 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n259), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n269), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n258), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n257), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n260) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_U60 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n285), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n264), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n256), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n257) );
  NAND4_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_U59 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n261), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n255), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n283), .A4(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n269), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n258) );
  AOI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_U58 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n278), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n254), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n253), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n284), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n259) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_U57 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n265), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n266), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n252), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n284) );
  NOR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_U56 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n285), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n251), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n287), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n253) );
  AND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_U55 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n265), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n266), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n287) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_U54 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n250), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n266) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_U53 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n256), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n276), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n278) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_U52 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n252), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n267), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n247), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n248) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_U51 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n250), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n246), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n264), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n247) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_U50 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n283), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n286), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n264) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_U49 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n269), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n276), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n286) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_U48 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n251), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n263), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n252) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_U47 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n245), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n254), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n263) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_U46 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n244), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n249) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_U45 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n276), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n255), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n268), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n244) );
  AND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_U44 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n250), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n246), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n268) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_U43 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n285), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n279), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n246) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_U42 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n256), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n280), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n250) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_U41 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n262), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n280) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_U40 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n256), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n254), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n255) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_U39 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n282), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n262), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n261) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_U38 ( .A(
        Red_StateRegOutput[60]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n243), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n262) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_U37 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n285), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n282) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_U36 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n276), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n251) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_U35 ( .A(
        Red_StateRegOutput[61]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n242), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n276) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_U34 ( .A(
        F_SD2_RedSB_inst_n50), .B(F_SD2_RedSB_inst_n52), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n242) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_U33 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n269), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n245), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n277) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_U32 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n256), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n245) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_U31 ( .A(
        Red_StateRegOutput[59]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n241), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n256) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_U30 ( .A(
        F_SD2_RedSB_inst_n49), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n240), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n269) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_U29 ( .A(
        Red_StateRegOutput[58]), .B(F_SD2_RedSB_inst_n51), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n240) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_U28 ( .A(
        F_SD2_RedSB_inst_n50), .B(F_SD2_RedSB_inst_n51), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n243) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_U27 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n283), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n254), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n265) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_U26 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n279), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n254) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_U25 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n239), .B(
        Red_StateRegOutput[62]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n279) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_U24 ( .A(
        F_SD2_RedSB_inst_n51), .B(F_SD2_RedSB_inst_n52), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n239) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_U23 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n267), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n283) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_U22 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n238), .B(
        Red_StateRegOutput[57]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n267) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_U21 ( .A(
        F_SD2_RedSB_inst_n50), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n241), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n238) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_U20 ( .A(
        F_SD2_RedSB_inst_n49), .B(F_SD2_RedSB_inst_n52), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n241) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_U19 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n235), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n234), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n236), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n237), .ZN(Red_Feedback[31])
         );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_U18 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n235), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n230), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n234), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n237) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_U17 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n289), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n290), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n291), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n236) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_U16 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n289), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n290), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n288), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n235) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_U15 ( .A(
        Red_StateRegOutput[57]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n233), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n234) );
  AOI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_U14 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n267), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n249), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n232), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n248), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n233) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_U13 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n265), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n231), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n232) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_U12 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n261), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n251), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n277), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n285), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n231) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_U11 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n291), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n230) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_U10 ( .A(
        Red_StateRegOutput[56]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n229), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n285) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_U9 ( .A(
        F_SD2_RedSB_inst_n49), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n243), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n229) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_U8 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n228), .B(
        Red_StateRegOutput[56]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n291) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_U7 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n224), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n284), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n227), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n228) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_U6 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n283), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n225), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n282), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n226), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n227) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_U5 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n281), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n279), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n280), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n226) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_U4 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n276), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n277), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n280), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n278), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n225) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_U3 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n287), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n286), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n285), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_59_n224) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_U73 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n277), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n276), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n279), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n278) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_U72 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n275), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n274), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n273), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n277) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_U71 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n272), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n279) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_U70 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n267), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n266), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n265), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n268) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_U69 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n263), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n262), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n280) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_U68 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n265), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n281), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n261), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n276) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_U67 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n265), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n260), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n283) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_U66 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n263), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n264), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n258), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n285), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n259) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_U65 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n272), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n257), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n285) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_U64 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n270), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n256), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n282) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_U63 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n286), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n274) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_U62 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n260), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n255), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n286) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_U61 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n262), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n271), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n254), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n252) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_U60 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n273), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n251), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n250), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n253) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_U59 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n284), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n250) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_U58 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n270), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n256), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n284) );
  OR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_U57 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n275), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n257), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n256) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_U56 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n267), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n270) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_U55 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n258), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n275), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n251) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_U54 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n281), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n258) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_U53 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n272), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n248), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n247), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n249) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_U52 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n262), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n264), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n246), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n245), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n247) );
  OR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_U51 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n254), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n271), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n269), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n245) );
  OR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_U50 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n281), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n257), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n263), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n269) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_U49 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n260), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n254) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_U48 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n267), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n255), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n266), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n244), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n257), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n246) );
  AND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_U47 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n267), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n255), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n244) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_U46 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n275), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n260), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n266) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_U45 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n265), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n281), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n255) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_U44 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n263), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n265) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_U43 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n272), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n273), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n267) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_U42 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n273), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n257), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n264) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_U41 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n271), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n273) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_U40 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n275), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n281), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n262) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_U39 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n261), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n275) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_U38 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n261), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n243), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n263), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n243), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n257), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n248) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_U37 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n242), .B(
        Red_StateRegOutput[56]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n257) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_U36 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n241), .B(
        F_SD2_RedSB_inst_n50), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n242) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_U35 ( .A(
        Red_StateRegOutput[58]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n241), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n263) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_U34 ( .A(
        F_SD2_RedSB_inst_n51), .B(F_SD2_RedSB_inst_n49), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n241) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_U33 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n260), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n281), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n271), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n243) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_U32 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n240), .B(
        Red_StateRegOutput[59]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n271) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_U31 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n239), .B(
        F_SD2_RedSB_inst_n50), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n281) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_U30 ( .A(
        Red_StateRegOutput[61]), .B(F_SD2_RedSB_inst_n52), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n239) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_U29 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n238), .B(
        Red_StateRegOutput[57]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n260) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_U28 ( .A(
        F_SD2_RedSB_inst_n50), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n240), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n238) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_U27 ( .A(
        F_SD2_RedSB_inst_n49), .B(F_SD2_RedSB_inst_n52), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n240) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_U26 ( .A(
        Red_StateRegOutput[62]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n237), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n261) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_U25 ( .A(
        F_SD2_RedSB_inst_n51), .B(F_SD2_RedSB_inst_n52), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n237) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_U24 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n236), .B(
        Red_StateRegOutput[60]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n272) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_U23 ( .A(
        F_SD2_RedSB_inst_n51), .B(F_SD2_RedSB_inst_n50), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n236) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_U22 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n217), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n221), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n234), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n225), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n235), .ZN(Red_Feedback[32])
         );
  NOR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_U21 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n221), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n225), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n234), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n235) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_U20 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n232), .B2(
        Red_StateRegOutput[58]), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n233), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n234) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_U19 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n232), .B2(
        Red_StateRegOutput[58]), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n217), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n233) );
  AOI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_U18 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n271), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n227), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n229), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n231), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n232) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_U17 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n271), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n230), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n264), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n286), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n231) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_U16 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n280), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n230) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_U15 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n270), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n228), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n268), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n269), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n229) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_U14 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n266), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n228) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_U13 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n285), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n226), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n276), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n227) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_U12 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n275), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n283), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n226) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_U11 ( .A(
        Red_StateRegOutput[61]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n224), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n225) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_U10 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n285), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n286), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n222), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n223), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n224) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_U9 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n279), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n280), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n278), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n223) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_U8 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n284), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n282), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n284), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n283), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n281), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n222) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_U7 ( .A(
        Red_StateRegOutput[57]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n220), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n221) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_U6 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n219), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n218), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n220) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_U5 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n254), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n253), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n252), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n219) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_U4 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n266), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n259), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n282), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n274), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n218) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_U3 ( .A(
        Red_StateRegOutput[56]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n249), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_60_n217) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_U73 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n284), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n283), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n282), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n281), .ZN(Red_Feedback[33])
         );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_U72 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n280), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n281), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n279), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n283) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_U71 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n280), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n281), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n282), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n279) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_U70 ( .A(
        Red_StateRegOutput[61]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n278), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n282) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_U69 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n277), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n276), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n278) );
  NAND4_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_U68 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n275), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n274), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n273), .A4(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n272), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n276) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_U67 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n271), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n270), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n269), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n268), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n277) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_U66 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n267), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n268) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_U65 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n274), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n266), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n265), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n264), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n270) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_U64 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n263), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n265) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_U63 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n262), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n272), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n261), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n260), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n266) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_U62 ( .A(
        Red_StateRegOutput[57]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n259), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n281) );
  NOR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_U61 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n258), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n257), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n256), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n259) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_U60 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n255), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n254), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n255), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n253), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n252), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n256) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_U59 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n273), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n263), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n252) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_U58 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n251), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n250), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n263) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_U57 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n275), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n262), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n253) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_U56 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n271), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n269), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n254) );
  AOI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_U55 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n275), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n249), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n248), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n247), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n257) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_U54 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n246), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n245), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n275), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n247) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_U53 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n271), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n244), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n249) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_U52 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n245), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n271) );
  NOR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_U51 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n251), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n244), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n250), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n258) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_U50 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n260), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n248), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n250) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_U49 ( .A(
        Red_StateRegOutput[56]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n243), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n280) );
  AOI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_U48 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n275), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n242), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n241), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n240), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n243) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_U47 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n251), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n239), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n255), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n238), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n240) );
  OR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_U46 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n251), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n239), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n260), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n238) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_U45 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n237), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n248), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n244), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n255) );
  NOR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_U44 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n237), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n236), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n272), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n241) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_U43 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n274), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n262), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n246), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n235), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n236) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_U42 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n234), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n260), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n233), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n242) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_U41 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n232), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n246), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n262), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n233) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_U40 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n231), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n234) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_U39 ( .A(
        Red_StateRegOutput[58]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n230), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n284) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_U38 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n262), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n229), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n228), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n230) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_U37 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n267), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n227), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n226), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n264), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n228) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_U36 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n244), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n225), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n264) );
  NAND4_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_U35 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n237), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n269), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n274), .A4(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n227), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n226) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_U34 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n272), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n269) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_U33 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n237), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n273), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n262), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n231), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n267) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_U32 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n245), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n248), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n231) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_U31 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n244), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n239), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n273) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_U30 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n245), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n225), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n239) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_U29 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n260), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n237) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_U28 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n274), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n224), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n223), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n251), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n229) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_U27 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n232), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n244), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n261), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n244), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n235), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n224) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_U26 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n275), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n245), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n235) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_U25 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n227), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n275) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_U24 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n251), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n261) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_U23 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n227), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n272), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n251) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_U22 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n222), .B(
        Red_StateRegOutput[60]), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n272) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_U21 ( .A(
        F_SD2_RedSB_inst_n50), .B(F_SD2_RedSB_inst_n51), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n222) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_U20 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n221), .B(
        Red_StateRegOutput[59]), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n227) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_U19 ( .A(
        F_SD2_RedSB_inst_n49), .B(F_SD2_RedSB_inst_n52), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n221) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_U18 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n246), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n244) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_U17 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n220), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n219), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n246) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_U16 ( .A(
        F_SD2_RedSB_inst_n52), .B(Red_StateRegOutput[57]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n220) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_U15 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n223), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n232) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_U14 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n260), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n245), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n223) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_U13 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n218), .B(
        Red_StateRegOutput[61]), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n245) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_U12 ( .A(
        F_SD2_RedSB_inst_n50), .B(F_SD2_RedSB_inst_n52), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n218) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_U11 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n217), .B(
        F_SD2_RedSB_inst_n51), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n260) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_U10 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n219), .B(
        Red_StateRegOutput[56]), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n217) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_U9 ( .A(
        F_SD2_RedSB_inst_n49), .B(F_SD2_RedSB_inst_n50), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n219) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_U8 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n248), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n274) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_U7 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n216), .B(
        Red_StateRegOutput[62]), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n248) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_U6 ( .A(
        F_SD2_RedSB_inst_n51), .B(F_SD2_RedSB_inst_n52), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n216) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_U5 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n225), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n262) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_U4 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n215), .B(
        F_SD2_RedSB_inst_n51), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n225) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_U3 ( .A(
        Red_StateRegOutput[58]), .B(F_SD2_RedSB_inst_n49), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_61_n215) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_U65 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n283), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n282), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n281), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n280), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n279), .ZN(Red_Feedback[34])
         );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_U64 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n283), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n282), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n281), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n279) );
  MUX2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_U63 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n283), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n282), .S(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n278), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n280) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_U62 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n277), .B(
        Red_StateRegOutput[58]), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n278) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_U61 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n276), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n275), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n274), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n277) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_U60 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n273), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n274) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_U59 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n272), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n271), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n270), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n269), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n268), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n273) );
  AND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_U58 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n267), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n266), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n265), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n269) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_U57 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n266), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n264), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n263), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n262), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n275) );
  AOI222_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_U56 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n261), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n260), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n261), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n259), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n260), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n259), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n263) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_U55 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n258), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n268), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n259) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_U54 ( .A(
        Red_StateRegOutput[56]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n257), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n281) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_U53 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n268), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n256), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n255), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n257) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_U52 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n268), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n254), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n262), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n255) );
  AOI222_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_U51 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n261), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n260), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n261), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n253), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n260), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n253), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n254) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_U50 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n276), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n258), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n253) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_U49 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n252), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n251), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n250), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n249), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n256) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_U48 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n276), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n266), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n248), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n247), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n252) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_U47 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n264), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n247) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_U46 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n272), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n258), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n264) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_U45 ( .A(
        Red_StateRegOutput[57]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n246), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n282) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_U44 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n248), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n262), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n245), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n244), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n246) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_U43 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n248), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n243), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n244) );
  AOI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_U42 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n271), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n242), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n241), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n240), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n245) );
  NOR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_U41 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n270), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n239), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n250), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n240) );
  AND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_U40 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n238), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n268), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n260), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n241) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_U39 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n248), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n266), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n260) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_U38 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n251), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n237), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n249), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n238) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_U37 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n276), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n270), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n249) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_U36 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n258), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n236), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n262) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_U35 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n237), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n258) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_U34 ( .A(
        Red_StateRegOutput[61]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n235), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n283) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_U33 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n234), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n237), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n233), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n237), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n232), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n235) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_U32 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n251), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n268), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n267), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n236), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n271), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n232) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_U31 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n250), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n276), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n271) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_U30 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n237), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n248), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n250) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_U29 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n239), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n272), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n236) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_U28 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n242), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n265), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n243), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n233) );
  AND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_U27 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n261), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n231), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n243) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_U26 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n276), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n248), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n265) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_U25 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n230), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n229), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n248) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_U24 ( .A(
        F_SD2_RedSB_inst_n49), .B(Red_StateRegOutput[57]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n230) );
  OR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_U23 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n261), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n231), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n242) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_U22 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n268), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n266), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n231) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_U21 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n228), .B(
        Red_StateRegOutput[56]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n268) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_U20 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n227), .B(
        F_SD2_RedSB_inst_n50), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n228) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_U19 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n267), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n270), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n261) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_U18 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n272), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n270) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_U17 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n226), .B(
        Red_StateRegOutput[59]), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n272) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_U16 ( .A(
        F_SD2_RedSB_inst_n49), .B(F_SD2_RedSB_inst_n52), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n226) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_U15 ( .A(
        Red_StateRegOutput[61]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n229), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n237) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_U14 ( .A(
        F_SD2_RedSB_inst_n52), .B(F_SD2_RedSB_inst_n50), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n229) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_U13 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n225), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n234) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_U12 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n267), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n239), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n224), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n225) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_U11 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n267), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n239), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n276), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n224) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_U10 ( .A(
        Red_StateRegOutput[58]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n227), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n276) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_U9 ( .A(
        F_SD2_RedSB_inst_n51), .B(F_SD2_RedSB_inst_n49), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n227) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_U8 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n266), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n239) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_U7 ( .A(
        Red_StateRegOutput[62]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n223), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n266) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_U6 ( .A(
        F_SD2_RedSB_inst_n51), .B(F_SD2_RedSB_inst_n52), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n223) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_U5 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n251), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n267) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_U4 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n222), .B(
        Red_StateRegOutput[60]), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n251) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_U3 ( .A(
        F_SD2_RedSB_inst_n51), .B(F_SD2_RedSB_inst_n50), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_62_n222) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_U69 ( .A(
        Red_StateRegOutput[64]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n280), .Z(Red_Feedback[49])
         );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_U68 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n279), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n278), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n280) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_U67 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n277), .B2(
        Red_StateRegOutput[65]), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n276), .C2(
        Red_StateRegOutput[68]), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n275), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n278) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_U66 ( .A1(
        Red_StateRegOutput[65]), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n277), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n276), .B2(
        Red_StateRegOutput[68]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n275) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_U65 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n274), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n273), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n276) );
  AOI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_U64 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n272), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n271), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n270), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n269), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n273) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_U63 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n268), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n267), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n266), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n265), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n264), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n269) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_U62 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n268), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n263), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n262), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n270) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_U61 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n268), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n263), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n261), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n262) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_U60 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n260), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n259), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n258), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n271) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_U59 ( .A(
        Red_StateRegOutput[63]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n257), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n274) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_U58 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n256), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n255), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n254), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n257) );
  OR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_U57 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n267), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n253), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n252), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n254) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_U56 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n251), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n250), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n249), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n252) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_U55 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n250), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n251), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n248), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n253) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_U54 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n247), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n246), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n245), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n244), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n255) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_U53 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n243), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n242), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n241), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n240), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n247) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_U52 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n239), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n238), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n240), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n237), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n236), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n277) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_U51 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n235), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n234), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n233), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n236) );
  AOI222_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_U50 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n251), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n249), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n251), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n232), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n249), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n232), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n234) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_U49 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n242), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n267), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n232) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_U48 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n263), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n246), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n249) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_U47 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n231), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n251) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_U46 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n256), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n230), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n237) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_U45 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n261), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n263), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n229), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n238) );
  NOR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_U44 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n267), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n244), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n259), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n229) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_U43 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n245), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n246), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n259) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_U42 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n268), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n228), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n244) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_U41 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n256), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n267) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_U40 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n242), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n245), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n261) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_U39 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n264), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n260), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n227), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n279) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_U38 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n246), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n226), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n225), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n227) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_U37 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n246), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n224), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n248), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n225) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_U36 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n235), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n248) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_U35 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n242), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n265), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n235) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_U34 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n239), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n228), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n265) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_U33 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n241), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n243), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n256), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n263), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n224) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_U32 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n240), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n245), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n243) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_U31 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n266), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n242), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n241) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_U30 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n272), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n223), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n258), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n226) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_U29 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n231), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n222), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n258) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_U28 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n240), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n228), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n223) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_U27 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n231), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n222), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n260) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_U26 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n228), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n256), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n222) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_U25 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n221), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n220), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n256) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_U24 ( .A(
        Red_StateRegOutput[63]), .B(F_SD2_RedSB_inst_n53), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n221) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_U23 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n263), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n228) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_U22 ( .A(
        Red_StateRegOutput[69]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n219), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n263) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_U21 ( .A(
        F_SD2_RedSB_inst_n56), .B(F_SD2_RedSB_inst_n55), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n219) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_U20 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n239), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n268), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n231) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_U19 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n266), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n268) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_U18 ( .A(
        Red_StateRegOutput[67]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n220), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n266) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_U17 ( .A(
        F_SD2_RedSB_inst_n54), .B(F_SD2_RedSB_inst_n55), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n220) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_U16 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n240), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n239) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_U15 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n218), .B(
        Red_StateRegOutput[66]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n240) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_U14 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n230), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n264) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_U13 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n250), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n246), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n230) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_U12 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n217), .B(
        F_SD2_RedSB_inst_n54), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n246) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_U11 ( .A(
        Red_StateRegOutput[64]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n218), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n217) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_U10 ( .A(
        F_SD2_RedSB_inst_n56), .B(F_SD2_RedSB_inst_n53), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n218) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_U9 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n242), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n245), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n250) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_U8 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n233), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n245) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_U7 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n216), .B(
        Red_StateRegOutput[65]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n233) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_U6 ( .A(
        F_SD2_RedSB_inst_n53), .B(F_SD2_RedSB_inst_n55), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n216) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_U5 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n272), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n242) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_U4 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n215), .B(
        F_SD2_RedSB_inst_n54), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n272) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_U3 ( .A(
        Red_StateRegOutput[68]), .B(F_SD2_RedSB_inst_n56), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_63_n215) );
  AOI222_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_U69 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n279), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n278), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n279), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n277), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n278), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n276), .ZN(Red_Feedback[50])
         );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_U68 ( .A(
        Red_StateRegOutput[68]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n275), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n276) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_U67 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n274), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n273), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n272), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n273), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n271), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n275) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_U66 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n270), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n269), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n268), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n269), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n267), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n271) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_U65 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n266), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n267) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_U64 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n265), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n264), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n268) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_U63 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n263), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n262), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n261), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n272) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_U62 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n260), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n259), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n262) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_U61 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n265), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n264), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n258), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n274) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_U60 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n265), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n264), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n257), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n258) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_U59 ( .A(
        Red_StateRegOutput[64]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n256), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n277) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_U58 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n255), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n254), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n253), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n256) );
  AOI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_U57 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n266), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n252), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n251), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n250), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n253) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_U56 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n249), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n248), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n260), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n261), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n250) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_U55 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n247), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n246), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n261) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_U54 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n245), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n260), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n244), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n243), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n249) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_U53 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n242), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n260) );
  NOR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_U52 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n241), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n240), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n239), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n251) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_U51 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n263), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n252) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_U50 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n247), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n246), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n263) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_U49 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n265), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n238), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n246) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_U48 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n244), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n238), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n254) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_U47 ( .A(
        Red_StateRegOutput[63]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n237), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n278) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_U46 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n238), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n236), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n235), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n237) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_U45 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n238), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n234), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n233), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n235) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_U44 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n244), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n247), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n259), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n248), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n233) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_U43 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n232), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n264), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n239), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n255), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n236) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_U42 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n257), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n241), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n255) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_U41 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n257), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n265), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n242), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n231), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n232) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_U40 ( .A(
        Red_StateRegOutput[65]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n230), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n279) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_U39 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n229), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n259), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n228), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n257), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n227), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n230) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_U38 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n226), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n225), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n224), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n223), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n227) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_U37 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n257), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n244), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n223) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_U36 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n222), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n224) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_U35 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n241), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n266), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n225) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_U34 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n257), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n239), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n266) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_U33 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n242), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n248), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n239) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_U32 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n259), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n257) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_U31 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n234), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n221), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n228) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_U30 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n222), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n247), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n231), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n240), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n221) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_U29 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n241), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n248), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n231) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_U28 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n273), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n248) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_U27 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n273), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n238), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n222) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_U26 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n273), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n245), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n244), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n247), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n234) );
  AND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_U25 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n270), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n264), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n247) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_U24 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n265), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n242), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n244) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_U23 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n240), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n265) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_U22 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n240), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n270), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n245) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_U21 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n241), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n270) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_U20 ( .A(
        Red_StateRegOutput[68]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n220), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n273) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_U19 ( .A(
        F_SD2_RedSB_inst_n55), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n219), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n259) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_U18 ( .A(
        Red_StateRegOutput[65]), .B(F_SD2_RedSB_inst_n53), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n219) );
  NOR4_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_U17 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n242), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n241), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n240), .A4(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n269), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n229) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_U16 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n243), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n269) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_U15 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n264), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n226), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n243) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_U14 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n238), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n226) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_U13 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n218), .B(
        Red_StateRegOutput[63]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n238) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_U12 ( .A(
        F_SD2_RedSB_inst_n53), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n217), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n218) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_U11 ( .A(
        Red_StateRegOutput[67]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n217), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n264) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_U10 ( .A(
        F_SD2_RedSB_inst_n55), .B(F_SD2_RedSB_inst_n54), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n217) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_U9 ( .A(
        Red_StateRegOutput[69]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n216), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n240) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_U8 ( .A(
        F_SD2_RedSB_inst_n55), .B(F_SD2_RedSB_inst_n56), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n216) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_U7 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n215), .B(
        Red_StateRegOutput[66]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n241) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_U6 ( .A(
        F_SD2_RedSB_inst_n53), .B(F_SD2_RedSB_inst_n56), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n215) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_U5 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n214), .B(
        Red_StateRegOutput[64]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n242) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_U4 ( .A(
        F_SD2_RedSB_inst_n53), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n220), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n214) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_U3 ( .A(
        F_SD2_RedSB_inst_n54), .B(F_SD2_RedSB_inst_n56), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_64_n220) );
  MUX2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_U54 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n240), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n239), .S(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n238), .Z(Red_Feedback[51])
         );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_U53 ( .A(
        Red_StateRegOutput[65]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n237), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n238) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_U52 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n236), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n235), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n234), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n233), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n237) );
  OR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_U51 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n232), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n231), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n230), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n233) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_U50 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n229), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n228), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n227), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n234) );
  AOI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_U49 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n226), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n225), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n224), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n223), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n236) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_U48 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n222), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n221), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n220), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n221), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n219), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n223) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_U47 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n226), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n225), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n218), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n221) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_U46 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n217), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n216), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n225) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_U45 ( .A(
        Red_StateRegOutput[68]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n215), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n239) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_U44 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n214), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n230), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n213), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n212), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n215) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_U43 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n228), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n226), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n211), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n232), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n212) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_U42 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n210), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n228), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n210), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n226), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n216), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n213) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_U41 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n220), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n216) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_U40 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n209), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n226) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_U39 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n208), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n207), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n228) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_U38 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n219), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n206), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n205), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n210) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_U37 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n219), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n206), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n208), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n205) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_U36 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n235), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n208) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_U35 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n222), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n204), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n229), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n214) );
  AND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_U34 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n206), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n219), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n204) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_U33 ( .A(
        Red_StateRegOutput[64]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n203), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n240) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_U32 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n202), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n201), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n200), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n201), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n199), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n203) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_U31 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n198), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n197), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n230), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n209), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n199) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_U30 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n227), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n220), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n218), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n197) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_U29 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n207), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n218) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_U28 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n222), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n201), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n227) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_U27 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n198), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n230), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n209), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n230), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n217), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n200) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_U26 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n231), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n206), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n209) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_U25 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n207), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n235), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n220), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n230) );
  AOI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_U24 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n229), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n211), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n207), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n224), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n198) );
  NOR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_U23 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n231), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n220), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n201), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n224) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_U22 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n219), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n220), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n211) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_U21 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n196), .B(
        Red_StateRegOutput[68]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n220) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_U20 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n201), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n219) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_U19 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n232), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n206), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n229) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_U18 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n195), .B(
        Red_StateRegOutput[67]), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n206) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_U17 ( .A(
        F_SD2_RedSB_inst_n55), .B(F_SD2_RedSB_inst_n54), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n195) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_U16 ( .A(
        Red_StateRegOutput[69]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n194), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n201) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_U15 ( .A(
        F_SD2_RedSB_inst_n55), .B(F_SD2_RedSB_inst_n56), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n194) );
  NOR4_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_U14 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n207), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n231), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n232), .A4(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n235), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n202) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_U13 ( .A(
        Red_StateRegOutput[65]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n193), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n235) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_U12 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n217), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n232) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_U11 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n192), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n193), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n217) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_U10 ( .A(
        F_SD2_RedSB_inst_n53), .B(F_SD2_RedSB_inst_n55), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n193) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_U9 ( .A(
        F_SD2_RedSB_inst_n54), .B(Red_StateRegOutput[63]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n192) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_U8 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n222), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n231) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_U7 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n191), .B(
        Red_StateRegOutput[66]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n222) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_U6 ( .A(
        F_SD2_RedSB_inst_n53), .B(F_SD2_RedSB_inst_n56), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n191) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_U5 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n190), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n196), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n207) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_U4 ( .A(
        F_SD2_RedSB_inst_n54), .B(F_SD2_RedSB_inst_n56), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n196) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_U3 ( .A(
        F_SD2_RedSB_inst_n53), .B(Red_StateRegOutput[64]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_65_n190) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_U71 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n289), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n291), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n290), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n288) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_U70 ( .A(
        Red_StateRegOutput[68]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n275), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n289) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_U69 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n274), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n273), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n272), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n276), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n275) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_U68 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n271), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n281), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n270), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n269), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n268), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n272) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_U67 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n267), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n266), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n285), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n265), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n270) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_U66 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n269), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n281) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_U65 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n280), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n279), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n271) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_U64 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n264), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n273) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_U63 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n263), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n262), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n261), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n274) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_U62 ( .A(
        Red_StateRegOutput[65]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n260), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n290) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_U61 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n259), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n269), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n258), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n257), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n260) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_U60 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n285), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n264), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n256), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n257) );
  NAND4_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_U59 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n261), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n255), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n283), .A4(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n269), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n258) );
  AOI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_U58 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n278), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n254), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n253), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n284), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n259) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_U57 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n265), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n266), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n252), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n284) );
  NOR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_U56 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n285), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n251), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n287), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n253) );
  AND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_U55 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n265), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n266), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n287) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_U54 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n250), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n266) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_U53 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n256), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n276), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n278) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_U52 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n252), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n267), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n247), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n248) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_U51 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n250), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n246), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n264), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n247) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_U50 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n283), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n286), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n264) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_U49 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n269), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n276), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n286) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_U48 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n251), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n263), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n252) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_U47 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n245), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n254), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n263) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_U46 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n244), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n249) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_U45 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n276), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n255), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n268), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n244) );
  AND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_U44 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n250), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n246), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n268) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_U43 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n285), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n279), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n246) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_U42 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n256), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n280), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n250) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_U41 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n262), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n280) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_U40 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n256), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n254), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n255) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_U39 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n282), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n262), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n261) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_U38 ( .A(
        Red_StateRegOutput[67]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n243), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n262) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_U37 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n285), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n282) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_U36 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n276), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n251) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_U35 ( .A(
        Red_StateRegOutput[68]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n242), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n276) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_U34 ( .A(
        F_SD2_RedSB_inst_n54), .B(F_SD2_RedSB_inst_n56), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n242) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_U33 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n269), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n245), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n277) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_U32 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n256), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n245) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_U31 ( .A(
        Red_StateRegOutput[66]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n241), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n256) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_U30 ( .A(
        F_SD2_RedSB_inst_n53), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n240), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n269) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_U29 ( .A(
        Red_StateRegOutput[65]), .B(F_SD2_RedSB_inst_n55), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n240) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_U28 ( .A(
        F_SD2_RedSB_inst_n54), .B(F_SD2_RedSB_inst_n55), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n243) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_U27 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n283), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n254), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n265) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_U26 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n279), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n254) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_U25 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n239), .B(
        Red_StateRegOutput[69]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n279) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_U24 ( .A(
        F_SD2_RedSB_inst_n55), .B(F_SD2_RedSB_inst_n56), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n239) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_U23 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n267), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n283) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_U22 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n238), .B(
        Red_StateRegOutput[64]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n267) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_U21 ( .A(
        F_SD2_RedSB_inst_n54), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n241), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n238) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_U20 ( .A(
        F_SD2_RedSB_inst_n53), .B(F_SD2_RedSB_inst_n56), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n241) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_U19 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n235), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n234), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n236), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n237), .ZN(Red_Feedback[52])
         );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_U18 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n235), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n230), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n234), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n237) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_U17 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n289), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n290), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n291), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n236) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_U16 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n289), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n290), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n288), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n235) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_U15 ( .A(
        Red_StateRegOutput[64]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n233), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n234) );
  AOI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_U14 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n267), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n249), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n232), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n248), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n233) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_U13 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n265), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n231), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n232) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_U12 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n261), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n251), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n277), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n285), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n231) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_U11 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n291), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n230) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_U10 ( .A(
        Red_StateRegOutput[63]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n229), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n285) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_U9 ( .A(
        F_SD2_RedSB_inst_n53), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n243), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n229) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_U8 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n228), .B(
        Red_StateRegOutput[63]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n291) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_U7 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n224), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n284), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n227), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n228) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_U6 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n283), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n225), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n282), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n226), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n227) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_U5 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n281), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n279), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n280), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n226) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_U4 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n276), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n277), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n280), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n278), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n225) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_U3 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n287), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n286), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n285), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_66_n224) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_U73 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n277), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n276), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n279), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n278) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_U72 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n275), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n274), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n273), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n277) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_U71 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n272), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n279) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_U70 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n267), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n266), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n265), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n268) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_U69 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n263), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n262), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n280) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_U68 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n265), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n281), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n261), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n276) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_U67 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n265), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n260), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n283) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_U66 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n263), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n264), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n258), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n285), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n259) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_U65 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n272), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n257), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n285) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_U64 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n270), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n256), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n282) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_U63 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n286), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n274) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_U62 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n260), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n255), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n286) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_U61 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n262), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n271), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n254), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n252) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_U60 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n273), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n251), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n250), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n253) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_U59 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n284), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n250) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_U58 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n270), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n256), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n284) );
  OR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_U57 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n275), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n257), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n256) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_U56 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n267), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n270) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_U55 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n258), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n275), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n251) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_U54 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n281), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n258) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_U53 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n272), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n248), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n247), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n249) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_U52 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n262), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n264), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n246), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n245), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n247) );
  OR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_U51 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n254), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n271), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n269), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n245) );
  OR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_U50 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n281), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n257), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n263), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n269) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_U49 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n260), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n254) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_U48 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n267), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n255), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n266), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n244), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n257), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n246) );
  AND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_U47 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n267), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n255), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n244) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_U46 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n275), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n260), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n266) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_U45 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n265), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n281), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n255) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_U44 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n263), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n265) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_U43 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n272), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n273), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n267) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_U42 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n273), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n257), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n264) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_U41 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n271), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n273) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_U40 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n275), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n281), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n262) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_U39 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n261), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n275) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_U38 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n261), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n243), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n263), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n243), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n257), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n248) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_U37 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n242), .B(
        Red_StateRegOutput[63]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n257) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_U36 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n241), .B(
        F_SD2_RedSB_inst_n54), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n242) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_U35 ( .A(
        Red_StateRegOutput[65]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n241), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n263) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_U34 ( .A(
        F_SD2_RedSB_inst_n55), .B(F_SD2_RedSB_inst_n53), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n241) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_U33 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n260), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n281), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n271), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n243) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_U32 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n240), .B(
        Red_StateRegOutput[66]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n271) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_U31 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n239), .B(
        F_SD2_RedSB_inst_n54), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n281) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_U30 ( .A(
        Red_StateRegOutput[68]), .B(F_SD2_RedSB_inst_n56), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n239) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_U29 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n238), .B(
        Red_StateRegOutput[64]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n260) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_U28 ( .A(
        F_SD2_RedSB_inst_n54), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n240), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n238) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_U27 ( .A(
        F_SD2_RedSB_inst_n53), .B(F_SD2_RedSB_inst_n56), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n240) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_U26 ( .A(
        Red_StateRegOutput[69]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n237), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n261) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_U25 ( .A(
        F_SD2_RedSB_inst_n55), .B(F_SD2_RedSB_inst_n56), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n237) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_U24 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n236), .B(
        Red_StateRegOutput[67]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n272) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_U23 ( .A(
        F_SD2_RedSB_inst_n55), .B(F_SD2_RedSB_inst_n54), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n236) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_U22 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n217), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n221), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n234), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n225), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n235), .ZN(Red_Feedback[53])
         );
  NOR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_U21 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n221), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n225), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n234), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n235) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_U20 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n232), .B2(
        Red_StateRegOutput[65]), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n233), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n234) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_U19 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n232), .B2(
        Red_StateRegOutput[65]), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n217), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n233) );
  AOI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_U18 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n271), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n227), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n229), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n231), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n232) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_U17 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n271), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n230), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n264), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n286), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n231) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_U16 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n280), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n230) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_U15 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n270), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n228), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n268), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n269), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n229) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_U14 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n266), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n228) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_U13 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n285), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n226), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n276), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n227) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_U12 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n275), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n283), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n226) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_U11 ( .A(
        Red_StateRegOutput[68]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n224), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n225) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_U10 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n285), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n286), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n222), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n223), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n224) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_U9 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n279), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n280), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n278), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n223) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_U8 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n284), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n282), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n284), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n283), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n281), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n222) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_U7 ( .A(
        Red_StateRegOutput[64]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n220), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n221) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_U6 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n219), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n218), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n220) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_U5 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n254), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n253), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n252), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n219) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_U4 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n266), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n259), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n282), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n274), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n218) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_U3 ( .A(
        Red_StateRegOutput[63]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n249), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_67_n217) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_U73 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n284), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n283), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n282), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n281), .ZN(Red_Feedback[54])
         );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_U72 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n280), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n281), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n279), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n283) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_U71 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n280), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n281), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n282), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n279) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_U70 ( .A(
        Red_StateRegOutput[68]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n278), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n282) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_U69 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n277), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n276), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n278) );
  NAND4_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_U68 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n275), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n274), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n273), .A4(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n272), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n276) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_U67 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n271), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n270), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n269), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n268), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n277) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_U66 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n267), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n268) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_U65 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n274), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n266), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n265), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n264), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n270) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_U64 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n263), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n265) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_U63 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n262), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n272), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n261), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n260), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n266) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_U62 ( .A(
        Red_StateRegOutput[64]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n259), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n281) );
  NOR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_U61 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n258), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n257), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n256), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n259) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_U60 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n255), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n254), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n255), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n253), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n252), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n256) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_U59 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n273), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n263), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n252) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_U58 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n251), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n250), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n263) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_U57 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n275), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n262), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n253) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_U56 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n271), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n269), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n254) );
  AOI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_U55 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n275), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n249), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n248), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n247), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n257) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_U54 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n246), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n245), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n275), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n247) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_U53 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n271), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n244), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n249) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_U52 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n245), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n271) );
  NOR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_U51 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n251), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n244), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n250), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n258) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_U50 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n260), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n248), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n250) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_U49 ( .A(
        Red_StateRegOutput[63]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n243), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n280) );
  AOI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_U48 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n275), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n242), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n241), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n240), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n243) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_U47 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n251), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n239), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n255), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n238), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n240) );
  OR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_U46 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n251), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n239), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n260), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n238) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_U45 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n237), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n248), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n244), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n255) );
  NOR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_U44 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n237), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n236), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n272), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n241) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_U43 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n274), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n262), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n246), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n235), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n236) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_U42 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n234), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n260), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n233), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n242) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_U41 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n232), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n246), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n262), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n233) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_U40 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n231), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n234) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_U39 ( .A(
        Red_StateRegOutput[65]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n230), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n284) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_U38 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n262), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n229), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n228), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n230) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_U37 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n267), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n227), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n226), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n264), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n228) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_U36 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n244), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n225), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n264) );
  NAND4_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_U35 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n237), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n269), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n274), .A4(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n227), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n226) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_U34 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n272), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n269) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_U33 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n237), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n273), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n262), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n231), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n267) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_U32 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n245), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n248), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n231) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_U31 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n244), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n239), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n273) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_U30 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n245), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n225), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n239) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_U29 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n260), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n237) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_U28 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n274), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n224), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n223), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n251), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n229) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_U27 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n232), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n244), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n261), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n244), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n235), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n224) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_U26 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n275), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n245), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n235) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_U25 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n227), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n275) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_U24 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n251), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n261) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_U23 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n227), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n272), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n251) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_U22 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n222), .B(
        Red_StateRegOutput[67]), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n272) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_U21 ( .A(
        F_SD2_RedSB_inst_n54), .B(F_SD2_RedSB_inst_n55), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n222) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_U20 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n221), .B(
        Red_StateRegOutput[66]), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n227) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_U19 ( .A(
        F_SD2_RedSB_inst_n53), .B(F_SD2_RedSB_inst_n56), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n221) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_U18 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n246), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n244) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_U17 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n220), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n219), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n246) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_U16 ( .A(
        F_SD2_RedSB_inst_n56), .B(Red_StateRegOutput[64]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n220) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_U15 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n223), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n232) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_U14 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n260), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n245), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n223) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_U13 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n218), .B(
        Red_StateRegOutput[68]), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n245) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_U12 ( .A(
        F_SD2_RedSB_inst_n54), .B(F_SD2_RedSB_inst_n56), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n218) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_U11 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n217), .B(
        F_SD2_RedSB_inst_n55), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n260) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_U10 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n219), .B(
        Red_StateRegOutput[63]), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n217) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_U9 ( .A(
        F_SD2_RedSB_inst_n53), .B(F_SD2_RedSB_inst_n54), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n219) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_U8 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n248), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n274) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_U7 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n216), .B(
        Red_StateRegOutput[69]), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n248) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_U6 ( .A(
        F_SD2_RedSB_inst_n55), .B(F_SD2_RedSB_inst_n56), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n216) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_U5 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n225), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n262) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_U4 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n215), .B(
        F_SD2_RedSB_inst_n55), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n225) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_U3 ( .A(
        Red_StateRegOutput[65]), .B(F_SD2_RedSB_inst_n53), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_68_n215) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_U65 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n283), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n282), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n281), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n280), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n279), .ZN(Red_Feedback[55])
         );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_U64 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n283), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n282), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n281), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n279) );
  MUX2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_U63 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n283), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n282), .S(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n278), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n280) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_U62 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n277), .B(
        Red_StateRegOutput[65]), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n278) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_U61 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n276), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n275), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n274), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n277) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_U60 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n273), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n274) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_U59 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n272), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n271), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n270), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n269), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n268), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n273) );
  AND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_U58 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n267), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n266), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n265), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n269) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_U57 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n266), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n264), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n263), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n262), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n275) );
  AOI222_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_U56 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n261), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n260), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n261), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n259), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n260), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n259), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n263) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_U55 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n258), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n268), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n259) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_U54 ( .A(
        Red_StateRegOutput[63]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n257), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n281) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_U53 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n268), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n256), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n255), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n257) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_U52 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n268), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n254), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n262), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n255) );
  AOI222_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_U51 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n261), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n260), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n261), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n253), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n260), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n253), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n254) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_U50 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n276), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n258), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n253) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_U49 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n252), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n251), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n250), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n249), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n256) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_U48 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n276), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n266), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n248), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n247), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n252) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_U47 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n264), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n247) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_U46 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n272), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n258), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n264) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_U45 ( .A(
        Red_StateRegOutput[64]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n246), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n282) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_U44 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n248), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n262), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n245), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n244), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n246) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_U43 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n248), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n243), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n244) );
  AOI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_U42 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n271), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n242), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n241), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n240), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n245) );
  NOR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_U41 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n270), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n239), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n250), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n240) );
  AND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_U40 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n238), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n268), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n260), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n241) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_U39 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n248), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n266), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n260) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_U38 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n251), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n237), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n249), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n238) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_U37 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n276), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n270), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n249) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_U36 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n258), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n236), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n262) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_U35 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n237), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n258) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_U34 ( .A(
        Red_StateRegOutput[68]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n235), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n283) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_U33 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n234), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n237), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n233), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n237), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n232), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n235) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_U32 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n251), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n268), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n267), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n236), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n271), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n232) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_U31 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n250), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n276), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n271) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_U30 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n237), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n248), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n250) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_U29 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n239), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n272), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n236) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_U28 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n242), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n265), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n243), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n233) );
  AND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_U27 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n261), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n231), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n243) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_U26 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n276), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n248), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n265) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_U25 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n230), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n229), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n248) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_U24 ( .A(
        F_SD2_RedSB_inst_n53), .B(Red_StateRegOutput[64]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n230) );
  OR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_U23 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n261), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n231), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n242) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_U22 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n268), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n266), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n231) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_U21 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n228), .B(
        Red_StateRegOutput[63]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n268) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_U20 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n227), .B(
        F_SD2_RedSB_inst_n54), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n228) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_U19 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n267), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n270), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n261) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_U18 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n272), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n270) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_U17 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n226), .B(
        Red_StateRegOutput[66]), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n272) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_U16 ( .A(
        F_SD2_RedSB_inst_n53), .B(F_SD2_RedSB_inst_n56), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n226) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_U15 ( .A(
        Red_StateRegOutput[68]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n229), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n237) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_U14 ( .A(
        F_SD2_RedSB_inst_n56), .B(F_SD2_RedSB_inst_n54), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n229) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_U13 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n225), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n234) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_U12 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n267), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n239), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n224), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n225) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_U11 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n267), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n239), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n276), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n224) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_U10 ( .A(
        Red_StateRegOutput[65]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n227), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n276) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_U9 ( .A(
        F_SD2_RedSB_inst_n55), .B(F_SD2_RedSB_inst_n53), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n227) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_U8 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n266), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n239) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_U7 ( .A(
        Red_StateRegOutput[69]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n223), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n266) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_U6 ( .A(
        F_SD2_RedSB_inst_n55), .B(F_SD2_RedSB_inst_n56), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n223) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_U5 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n251), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n267) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_U4 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n222), .B(
        Red_StateRegOutput[67]), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n251) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_U3 ( .A(
        F_SD2_RedSB_inst_n55), .B(F_SD2_RedSB_inst_n54), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_69_n222) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_U69 ( .A(
        Red_StateRegOutput[71]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n280), .Z(Red_Feedback[42])
         );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_U68 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n279), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n278), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n280) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_U67 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n277), .B2(
        Red_StateRegOutput[72]), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n276), .C2(
        Red_StateRegOutput[75]), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n275), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n278) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_U66 ( .A1(
        Red_StateRegOutput[72]), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n277), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n276), .B2(
        Red_StateRegOutput[75]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n275) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_U65 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n274), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n273), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n276) );
  AOI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_U64 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n272), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n271), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n270), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n269), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n273) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_U63 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n268), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n267), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n266), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n265), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n264), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n269) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_U62 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n268), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n263), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n262), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n270) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_U61 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n268), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n263), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n261), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n262) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_U60 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n260), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n259), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n258), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n271) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_U59 ( .A(
        Red_StateRegOutput[70]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n257), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n274) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_U58 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n256), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n255), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n254), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n257) );
  OR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_U57 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n267), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n253), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n252), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n254) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_U56 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n251), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n250), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n249), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n252) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_U55 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n250), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n251), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n248), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n253) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_U54 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n247), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n246), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n245), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n244), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n255) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_U53 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n243), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n242), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n241), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n240), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n247) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_U52 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n239), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n238), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n240), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n237), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n236), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n277) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_U51 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n235), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n234), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n233), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n236) );
  AOI222_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_U50 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n251), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n249), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n251), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n232), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n249), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n232), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n234) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_U49 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n242), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n267), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n232) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_U48 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n263), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n246), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n249) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_U47 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n231), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n251) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_U46 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n256), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n230), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n237) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_U45 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n261), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n263), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n229), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n238) );
  NOR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_U44 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n267), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n244), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n259), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n229) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_U43 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n245), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n246), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n259) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_U42 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n268), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n228), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n244) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_U41 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n256), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n267) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_U40 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n242), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n245), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n261) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_U39 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n264), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n260), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n227), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n279) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_U38 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n246), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n226), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n225), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n227) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_U37 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n246), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n224), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n248), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n225) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_U36 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n235), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n248) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_U35 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n242), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n265), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n235) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_U34 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n239), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n228), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n265) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_U33 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n241), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n243), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n256), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n263), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n224) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_U32 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n240), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n245), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n243) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_U31 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n266), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n242), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n241) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_U30 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n272), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n223), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n258), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n226) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_U29 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n231), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n222), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n258) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_U28 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n240), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n228), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n223) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_U27 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n231), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n222), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n260) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_U26 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n228), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n256), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n222) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_U25 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n221), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n220), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n256) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_U24 ( .A(
        Red_StateRegOutput[70]), .B(F_SD2_RedSB_inst_n57), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n221) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_U23 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n263), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n228) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_U22 ( .A(
        Red_StateRegOutput[76]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n219), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n263) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_U21 ( .A(
        F_SD2_RedSB_inst_n60), .B(F_SD2_RedSB_inst_n59), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n219) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_U20 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n239), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n268), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n231) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_U19 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n266), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n268) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_U18 ( .A(
        Red_StateRegOutput[74]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n220), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n266) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_U17 ( .A(
        F_SD2_RedSB_inst_n58), .B(F_SD2_RedSB_inst_n59), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n220) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_U16 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n240), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n239) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_U15 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n218), .B(
        Red_StateRegOutput[73]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n240) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_U14 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n230), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n264) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_U13 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n250), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n246), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n230) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_U12 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n217), .B(
        F_SD2_RedSB_inst_n58), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n246) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_U11 ( .A(
        Red_StateRegOutput[71]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n218), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n217) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_U10 ( .A(
        F_SD2_RedSB_inst_n60), .B(F_SD2_RedSB_inst_n57), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n218) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_U9 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n242), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n245), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n250) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_U8 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n233), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n245) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_U7 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n216), .B(
        Red_StateRegOutput[72]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n233) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_U6 ( .A(
        F_SD2_RedSB_inst_n57), .B(F_SD2_RedSB_inst_n59), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n216) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_U5 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n272), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n242) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_U4 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n215), .B(
        F_SD2_RedSB_inst_n58), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n272) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_U3 ( .A(
        Red_StateRegOutput[75]), .B(F_SD2_RedSB_inst_n60), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_70_n215) );
  AOI222_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_U69 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n279), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n278), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n279), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n277), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n278), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n276), .ZN(Red_Feedback[43])
         );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_U68 ( .A(
        Red_StateRegOutput[75]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n275), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n276) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_U67 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n274), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n273), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n272), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n273), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n271), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n275) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_U66 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n270), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n269), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n268), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n269), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n267), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n271) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_U65 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n266), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n267) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_U64 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n265), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n264), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n268) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_U63 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n263), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n262), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n261), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n272) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_U62 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n260), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n259), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n262) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_U61 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n265), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n264), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n258), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n274) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_U60 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n265), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n264), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n257), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n258) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_U59 ( .A(
        Red_StateRegOutput[71]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n256), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n277) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_U58 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n255), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n254), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n253), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n256) );
  AOI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_U57 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n266), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n252), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n251), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n250), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n253) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_U56 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n249), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n248), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n260), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n261), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n250) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_U55 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n247), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n246), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n261) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_U54 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n245), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n260), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n244), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n243), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n249) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_U53 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n242), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n260) );
  NOR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_U52 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n241), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n240), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n239), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n251) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_U51 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n263), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n252) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_U50 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n247), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n246), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n263) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_U49 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n265), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n238), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n246) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_U48 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n244), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n238), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n254) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_U47 ( .A(
        Red_StateRegOutput[70]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n237), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n278) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_U46 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n238), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n236), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n235), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n237) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_U45 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n238), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n234), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n233), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n235) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_U44 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n244), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n247), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n259), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n248), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n233) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_U43 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n232), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n264), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n239), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n255), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n236) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_U42 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n257), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n241), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n255) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_U41 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n257), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n265), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n242), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n231), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n232) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_U40 ( .A(
        Red_StateRegOutput[72]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n230), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n279) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_U39 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n229), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n259), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n228), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n257), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n227), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n230) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_U38 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n226), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n225), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n224), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n223), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n227) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_U37 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n257), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n244), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n223) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_U36 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n222), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n224) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_U35 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n241), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n266), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n225) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_U34 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n257), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n239), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n266) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_U33 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n242), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n248), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n239) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_U32 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n259), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n257) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_U31 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n234), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n221), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n228) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_U30 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n222), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n247), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n231), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n240), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n221) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_U29 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n241), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n248), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n231) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_U28 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n273), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n248) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_U27 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n273), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n238), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n222) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_U26 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n273), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n245), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n244), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n247), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n234) );
  AND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_U25 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n270), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n264), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n247) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_U24 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n265), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n242), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n244) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_U23 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n240), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n265) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_U22 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n240), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n270), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n245) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_U21 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n241), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n270) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_U20 ( .A(
        Red_StateRegOutput[75]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n220), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n273) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_U19 ( .A(
        F_SD2_RedSB_inst_n59), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n219), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n259) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_U18 ( .A(
        Red_StateRegOutput[72]), .B(F_SD2_RedSB_inst_n57), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n219) );
  NOR4_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_U17 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n242), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n241), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n240), .A4(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n269), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n229) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_U16 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n243), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n269) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_U15 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n264), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n226), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n243) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_U14 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n238), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n226) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_U13 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n218), .B(
        Red_StateRegOutput[70]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n238) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_U12 ( .A(
        F_SD2_RedSB_inst_n57), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n217), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n218) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_U11 ( .A(
        Red_StateRegOutput[74]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n217), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n264) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_U10 ( .A(
        F_SD2_RedSB_inst_n59), .B(F_SD2_RedSB_inst_n58), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n217) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_U9 ( .A(
        Red_StateRegOutput[76]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n216), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n240) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_U8 ( .A(
        F_SD2_RedSB_inst_n59), .B(F_SD2_RedSB_inst_n60), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n216) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_U7 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n215), .B(
        Red_StateRegOutput[73]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n241) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_U6 ( .A(
        F_SD2_RedSB_inst_n57), .B(F_SD2_RedSB_inst_n60), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n215) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_U5 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n214), .B(
        Red_StateRegOutput[71]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n242) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_U4 ( .A(
        F_SD2_RedSB_inst_n57), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n220), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n214) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_U3 ( .A(
        F_SD2_RedSB_inst_n58), .B(F_SD2_RedSB_inst_n60), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_71_n220) );
  MUX2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_U54 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n240), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n239), .S(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n238), .Z(Red_Feedback[44])
         );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_U53 ( .A(
        Red_StateRegOutput[72]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n237), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n238) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_U52 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n236), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n235), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n234), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n233), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n237) );
  OR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_U51 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n232), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n231), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n230), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n233) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_U50 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n229), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n228), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n227), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n234) );
  AOI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_U49 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n226), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n225), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n224), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n223), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n236) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_U48 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n222), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n221), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n220), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n221), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n219), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n223) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_U47 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n226), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n225), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n218), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n221) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_U46 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n217), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n216), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n225) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_U45 ( .A(
        Red_StateRegOutput[75]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n215), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n239) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_U44 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n214), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n230), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n213), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n212), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n215) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_U43 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n228), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n226), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n211), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n232), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n212) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_U42 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n210), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n228), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n210), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n226), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n216), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n213) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_U41 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n220), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n216) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_U40 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n209), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n226) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_U39 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n208), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n207), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n228) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_U38 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n219), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n206), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n205), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n210) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_U37 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n219), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n206), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n208), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n205) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_U36 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n235), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n208) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_U35 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n222), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n204), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n229), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n214) );
  AND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_U34 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n206), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n219), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n204) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_U33 ( .A(
        Red_StateRegOutput[71]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n203), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n240) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_U32 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n202), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n201), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n200), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n201), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n199), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n203) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_U31 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n198), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n197), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n230), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n209), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n199) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_U30 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n227), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n220), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n218), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n197) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_U29 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n207), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n218) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_U28 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n222), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n201), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n227) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_U27 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n198), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n230), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n209), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n230), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n217), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n200) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_U26 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n231), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n206), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n209) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_U25 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n207), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n235), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n220), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n230) );
  AOI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_U24 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n229), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n211), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n207), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n224), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n198) );
  NOR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_U23 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n231), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n220), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n201), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n224) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_U22 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n219), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n220), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n211) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_U21 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n196), .B(
        Red_StateRegOutput[75]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n220) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_U20 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n201), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n219) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_U19 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n232), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n206), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n229) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_U18 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n195), .B(
        Red_StateRegOutput[74]), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n206) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_U17 ( .A(
        F_SD2_RedSB_inst_n59), .B(F_SD2_RedSB_inst_n58), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n195) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_U16 ( .A(
        Red_StateRegOutput[76]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n194), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n201) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_U15 ( .A(
        F_SD2_RedSB_inst_n59), .B(F_SD2_RedSB_inst_n60), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n194) );
  NOR4_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_U14 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n207), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n231), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n232), .A4(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n235), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n202) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_U13 ( .A(
        Red_StateRegOutput[72]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n193), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n235) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_U12 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n217), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n232) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_U11 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n192), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n193), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n217) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_U10 ( .A(
        F_SD2_RedSB_inst_n57), .B(F_SD2_RedSB_inst_n59), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n193) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_U9 ( .A(
        F_SD2_RedSB_inst_n58), .B(Red_StateRegOutput[70]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n192) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_U8 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n222), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n231) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_U7 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n191), .B(
        Red_StateRegOutput[73]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n222) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_U6 ( .A(
        F_SD2_RedSB_inst_n57), .B(F_SD2_RedSB_inst_n60), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n191) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_U5 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n190), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n196), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n207) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_U4 ( .A(
        F_SD2_RedSB_inst_n58), .B(F_SD2_RedSB_inst_n60), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n196) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_U3 ( .A(
        F_SD2_RedSB_inst_n57), .B(Red_StateRegOutput[71]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_72_n190) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_U71 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n289), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n291), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n290), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n288) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_U70 ( .A(
        Red_StateRegOutput[75]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n275), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n289) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_U69 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n274), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n273), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n272), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n276), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n275) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_U68 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n271), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n281), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n270), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n269), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n268), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n272) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_U67 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n267), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n266), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n285), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n265), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n270) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_U66 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n269), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n281) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_U65 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n280), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n279), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n271) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_U64 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n264), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n273) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_U63 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n263), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n262), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n261), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n274) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_U62 ( .A(
        Red_StateRegOutput[72]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n260), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n290) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_U61 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n259), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n269), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n258), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n257), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n260) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_U60 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n285), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n264), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n256), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n257) );
  NAND4_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_U59 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n261), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n255), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n283), .A4(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n269), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n258) );
  AOI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_U58 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n278), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n254), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n253), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n284), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n259) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_U57 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n265), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n266), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n252), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n284) );
  NOR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_U56 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n285), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n251), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n287), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n253) );
  AND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_U55 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n265), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n266), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n287) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_U54 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n250), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n266) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_U53 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n256), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n276), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n278) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_U52 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n252), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n267), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n247), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n248) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_U51 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n250), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n246), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n264), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n247) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_U50 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n283), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n286), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n264) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_U49 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n269), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n276), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n286) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_U48 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n251), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n263), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n252) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_U47 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n245), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n254), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n263) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_U46 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n244), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n249) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_U45 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n276), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n255), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n268), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n244) );
  AND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_U44 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n250), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n246), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n268) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_U43 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n285), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n279), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n246) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_U42 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n256), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n280), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n250) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_U41 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n262), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n280) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_U40 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n256), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n254), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n255) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_U39 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n282), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n262), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n261) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_U38 ( .A(
        Red_StateRegOutput[74]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n243), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n262) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_U37 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n285), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n282) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_U36 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n276), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n251) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_U35 ( .A(
        Red_StateRegOutput[75]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n242), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n276) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_U34 ( .A(
        F_SD2_RedSB_inst_n58), .B(F_SD2_RedSB_inst_n60), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n242) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_U33 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n269), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n245), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n277) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_U32 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n256), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n245) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_U31 ( .A(
        Red_StateRegOutput[73]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n241), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n256) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_U30 ( .A(
        F_SD2_RedSB_inst_n57), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n240), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n269) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_U29 ( .A(
        Red_StateRegOutput[72]), .B(F_SD2_RedSB_inst_n59), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n240) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_U28 ( .A(
        F_SD2_RedSB_inst_n58), .B(F_SD2_RedSB_inst_n59), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n243) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_U27 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n283), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n254), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n265) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_U26 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n279), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n254) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_U25 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n239), .B(
        Red_StateRegOutput[76]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n279) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_U24 ( .A(
        F_SD2_RedSB_inst_n59), .B(F_SD2_RedSB_inst_n60), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n239) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_U23 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n267), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n283) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_U22 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n238), .B(
        Red_StateRegOutput[71]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n267) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_U21 ( .A(
        F_SD2_RedSB_inst_n58), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n241), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n238) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_U20 ( .A(
        F_SD2_RedSB_inst_n57), .B(F_SD2_RedSB_inst_n60), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n241) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_U19 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n235), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n234), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n236), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n237), .ZN(Red_Feedback[45])
         );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_U18 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n235), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n230), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n234), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n237) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_U17 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n289), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n290), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n291), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n236) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_U16 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n289), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n290), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n288), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n235) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_U15 ( .A(
        Red_StateRegOutput[71]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n233), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n234) );
  AOI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_U14 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n267), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n249), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n232), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n248), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n233) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_U13 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n265), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n231), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n232) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_U12 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n261), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n251), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n277), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n285), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n231) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_U11 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n291), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n230) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_U10 ( .A(
        Red_StateRegOutput[70]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n229), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n285) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_U9 ( .A(
        F_SD2_RedSB_inst_n57), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n243), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n229) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_U8 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n228), .B(
        Red_StateRegOutput[70]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n291) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_U7 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n224), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n284), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n227), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n228) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_U6 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n283), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n225), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n282), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n226), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n227) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_U5 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n281), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n279), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n280), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n226) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_U4 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n276), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n277), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n280), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n278), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n225) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_U3 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n287), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n286), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n285), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_73_n224) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_U73 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n277), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n276), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n279), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n278) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_U72 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n275), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n274), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n273), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n277) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_U71 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n272), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n279) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_U70 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n267), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n266), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n265), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n268) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_U69 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n263), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n262), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n280) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_U68 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n265), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n281), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n261), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n276) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_U67 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n265), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n260), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n283) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_U66 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n263), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n264), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n258), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n285), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n259) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_U65 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n272), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n257), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n285) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_U64 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n270), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n256), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n282) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_U63 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n286), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n274) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_U62 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n260), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n255), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n286) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_U61 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n262), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n271), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n254), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n252) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_U60 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n273), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n251), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n250), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n253) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_U59 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n284), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n250) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_U58 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n270), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n256), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n284) );
  OR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_U57 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n275), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n257), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n256) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_U56 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n267), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n270) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_U55 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n258), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n275), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n251) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_U54 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n281), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n258) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_U53 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n272), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n248), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n247), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n249) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_U52 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n262), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n264), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n246), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n245), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n247) );
  OR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_U51 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n254), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n271), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n269), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n245) );
  OR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_U50 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n281), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n257), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n263), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n269) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_U49 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n260), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n254) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_U48 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n267), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n255), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n266), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n244), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n257), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n246) );
  AND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_U47 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n267), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n255), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n244) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_U46 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n275), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n260), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n266) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_U45 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n265), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n281), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n255) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_U44 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n263), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n265) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_U43 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n272), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n273), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n267) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_U42 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n273), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n257), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n264) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_U41 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n271), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n273) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_U40 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n275), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n281), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n262) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_U39 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n261), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n275) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_U38 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n261), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n243), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n263), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n243), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n257), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n248) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_U37 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n242), .B(
        Red_StateRegOutput[70]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n257) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_U36 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n241), .B(
        F_SD2_RedSB_inst_n58), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n242) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_U35 ( .A(
        Red_StateRegOutput[72]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n241), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n263) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_U34 ( .A(
        F_SD2_RedSB_inst_n59), .B(F_SD2_RedSB_inst_n57), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n241) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_U33 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n260), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n281), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n271), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n243) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_U32 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n240), .B(
        Red_StateRegOutput[73]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n271) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_U31 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n239), .B(
        F_SD2_RedSB_inst_n58), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n281) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_U30 ( .A(
        Red_StateRegOutput[75]), .B(F_SD2_RedSB_inst_n60), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n239) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_U29 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n238), .B(
        Red_StateRegOutput[71]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n260) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_U28 ( .A(
        F_SD2_RedSB_inst_n58), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n240), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n238) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_U27 ( .A(
        F_SD2_RedSB_inst_n57), .B(F_SD2_RedSB_inst_n60), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n240) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_U26 ( .A(
        Red_StateRegOutput[76]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n237), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n261) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_U25 ( .A(
        F_SD2_RedSB_inst_n59), .B(F_SD2_RedSB_inst_n60), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n237) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_U24 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n236), .B(
        Red_StateRegOutput[74]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n272) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_U23 ( .A(
        F_SD2_RedSB_inst_n59), .B(F_SD2_RedSB_inst_n58), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n236) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_U22 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n217), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n221), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n234), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n225), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n235), .ZN(Red_Feedback[46])
         );
  NOR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_U21 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n221), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n225), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n234), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n235) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_U20 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n232), .B2(
        Red_StateRegOutput[72]), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n233), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n234) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_U19 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n232), .B2(
        Red_StateRegOutput[72]), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n217), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n233) );
  AOI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_U18 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n271), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n227), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n229), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n231), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n232) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_U17 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n271), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n230), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n264), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n286), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n231) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_U16 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n280), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n230) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_U15 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n270), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n228), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n268), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n269), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n229) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_U14 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n266), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n228) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_U13 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n285), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n226), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n276), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n227) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_U12 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n275), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n283), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n226) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_U11 ( .A(
        Red_StateRegOutput[75]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n224), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n225) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_U10 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n285), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n286), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n222), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n223), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n224) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_U9 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n279), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n280), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n278), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n223) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_U8 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n284), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n282), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n284), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n283), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n281), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n222) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_U7 ( .A(
        Red_StateRegOutput[71]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n220), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n221) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_U6 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n219), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n218), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n220) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_U5 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n254), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n253), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n252), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n219) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_U4 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n266), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n259), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n282), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n274), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n218) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_U3 ( .A(
        Red_StateRegOutput[70]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n249), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_74_n217) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_U73 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n284), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n283), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n282), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n281), .ZN(Red_Feedback[47])
         );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_U72 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n280), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n281), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n279), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n283) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_U71 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n280), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n281), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n282), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n279) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_U70 ( .A(
        Red_StateRegOutput[75]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n278), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n282) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_U69 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n277), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n276), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n278) );
  NAND4_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_U68 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n275), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n274), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n273), .A4(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n272), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n276) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_U67 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n271), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n270), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n269), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n268), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n277) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_U66 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n267), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n268) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_U65 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n274), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n266), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n265), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n264), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n270) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_U64 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n263), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n265) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_U63 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n262), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n272), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n261), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n260), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n266) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_U62 ( .A(
        Red_StateRegOutput[71]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n259), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n281) );
  NOR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_U61 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n258), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n257), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n256), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n259) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_U60 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n255), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n254), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n255), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n253), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n252), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n256) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_U59 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n273), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n263), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n252) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_U58 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n251), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n250), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n263) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_U57 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n275), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n262), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n253) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_U56 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n271), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n269), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n254) );
  AOI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_U55 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n275), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n249), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n248), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n247), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n257) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_U54 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n246), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n245), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n275), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n247) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_U53 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n271), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n244), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n249) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_U52 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n245), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n271) );
  NOR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_U51 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n251), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n244), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n250), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n258) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_U50 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n260), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n248), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n250) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_U49 ( .A(
        Red_StateRegOutput[70]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n243), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n280) );
  AOI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_U48 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n275), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n242), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n241), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n240), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n243) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_U47 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n251), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n239), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n255), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n238), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n240) );
  OR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_U46 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n251), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n239), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n260), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n238) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_U45 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n237), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n248), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n244), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n255) );
  NOR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_U44 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n237), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n236), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n272), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n241) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_U43 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n274), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n262), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n246), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n235), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n236) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_U42 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n234), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n260), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n233), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n242) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_U41 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n232), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n246), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n262), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n233) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_U40 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n231), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n234) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_U39 ( .A(
        Red_StateRegOutput[72]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n230), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n284) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_U38 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n262), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n229), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n228), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n230) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_U37 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n267), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n227), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n226), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n264), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n228) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_U36 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n244), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n225), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n264) );
  NAND4_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_U35 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n237), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n269), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n274), .A4(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n227), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n226) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_U34 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n272), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n269) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_U33 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n237), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n273), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n262), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n231), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n267) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_U32 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n245), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n248), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n231) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_U31 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n244), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n239), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n273) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_U30 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n245), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n225), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n239) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_U29 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n260), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n237) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_U28 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n274), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n224), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n223), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n251), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n229) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_U27 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n232), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n244), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n261), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n244), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n235), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n224) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_U26 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n275), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n245), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n235) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_U25 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n227), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n275) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_U24 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n251), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n261) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_U23 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n227), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n272), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n251) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_U22 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n222), .B(
        Red_StateRegOutput[74]), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n272) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_U21 ( .A(
        F_SD2_RedSB_inst_n58), .B(F_SD2_RedSB_inst_n59), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n222) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_U20 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n221), .B(
        Red_StateRegOutput[73]), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n227) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_U19 ( .A(
        F_SD2_RedSB_inst_n57), .B(F_SD2_RedSB_inst_n60), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n221) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_U18 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n246), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n244) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_U17 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n220), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n219), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n246) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_U16 ( .A(
        F_SD2_RedSB_inst_n60), .B(Red_StateRegOutput[71]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n220) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_U15 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n223), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n232) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_U14 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n260), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n245), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n223) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_U13 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n218), .B(
        Red_StateRegOutput[75]), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n245) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_U12 ( .A(
        F_SD2_RedSB_inst_n58), .B(F_SD2_RedSB_inst_n60), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n218) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_U11 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n217), .B(
        F_SD2_RedSB_inst_n59), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n260) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_U10 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n219), .B(
        Red_StateRegOutput[70]), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n217) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_U9 ( .A(
        F_SD2_RedSB_inst_n57), .B(F_SD2_RedSB_inst_n58), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n219) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_U8 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n248), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n274) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_U7 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n216), .B(
        Red_StateRegOutput[76]), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n248) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_U6 ( .A(
        F_SD2_RedSB_inst_n59), .B(F_SD2_RedSB_inst_n60), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n216) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_U5 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n225), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n262) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_U4 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n215), .B(
        F_SD2_RedSB_inst_n59), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n225) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_U3 ( .A(
        Red_StateRegOutput[72]), .B(F_SD2_RedSB_inst_n57), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_75_n215) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_U65 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n283), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n282), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n281), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n280), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n279), .ZN(Red_Feedback[48])
         );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_U64 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n283), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n282), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n281), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n279) );
  MUX2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_U63 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n283), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n282), .S(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n278), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n280) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_U62 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n277), .B(
        Red_StateRegOutput[72]), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n278) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_U61 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n276), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n275), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n274), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n277) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_U60 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n273), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n274) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_U59 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n272), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n271), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n270), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n269), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n268), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n273) );
  AND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_U58 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n267), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n266), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n265), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n269) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_U57 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n266), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n264), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n263), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n262), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n275) );
  AOI222_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_U56 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n261), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n260), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n261), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n259), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n260), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n259), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n263) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_U55 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n258), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n268), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n259) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_U54 ( .A(
        Red_StateRegOutput[70]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n257), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n281) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_U53 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n268), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n256), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n255), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n257) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_U52 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n268), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n254), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n262), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n255) );
  AOI222_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_U51 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n261), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n260), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n261), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n253), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n260), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n253), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n254) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_U50 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n276), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n258), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n253) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_U49 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n252), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n251), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n250), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n249), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n256) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_U48 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n276), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n266), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n248), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n247), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n252) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_U47 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n264), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n247) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_U46 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n272), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n258), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n264) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_U45 ( .A(
        Red_StateRegOutput[71]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n246), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n282) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_U44 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n248), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n262), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n245), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n244), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n246) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_U43 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n248), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n243), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n244) );
  AOI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_U42 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n271), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n242), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n241), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n240), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n245) );
  NOR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_U41 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n270), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n239), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n250), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n240) );
  AND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_U40 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n238), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n268), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n260), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n241) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_U39 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n248), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n266), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n260) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_U38 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n251), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n237), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n249), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n238) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_U37 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n276), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n270), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n249) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_U36 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n258), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n236), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n262) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_U35 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n237), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n258) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_U34 ( .A(
        Red_StateRegOutput[75]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n235), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n283) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_U33 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n234), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n237), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n233), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n237), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n232), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n235) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_U32 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n251), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n268), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n267), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n236), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n271), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n232) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_U31 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n250), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n276), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n271) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_U30 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n237), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n248), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n250) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_U29 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n239), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n272), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n236) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_U28 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n242), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n265), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n243), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n233) );
  AND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_U27 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n261), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n231), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n243) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_U26 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n276), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n248), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n265) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_U25 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n230), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n229), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n248) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_U24 ( .A(
        F_SD2_RedSB_inst_n57), .B(Red_StateRegOutput[71]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n230) );
  OR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_U23 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n261), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n231), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n242) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_U22 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n268), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n266), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n231) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_U21 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n228), .B(
        Red_StateRegOutput[70]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n268) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_U20 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n227), .B(
        F_SD2_RedSB_inst_n58), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n228) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_U19 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n267), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n270), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n261) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_U18 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n272), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n270) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_U17 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n226), .B(
        Red_StateRegOutput[73]), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n272) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_U16 ( .A(
        F_SD2_RedSB_inst_n57), .B(F_SD2_RedSB_inst_n60), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n226) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_U15 ( .A(
        Red_StateRegOutput[75]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n229), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n237) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_U14 ( .A(
        F_SD2_RedSB_inst_n60), .B(F_SD2_RedSB_inst_n58), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n229) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_U13 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n225), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n234) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_U12 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n267), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n239), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n224), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n225) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_U11 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n267), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n239), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n276), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n224) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_U10 ( .A(
        Red_StateRegOutput[72]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n227), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n276) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_U9 ( .A(
        F_SD2_RedSB_inst_n59), .B(F_SD2_RedSB_inst_n57), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n227) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_U8 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n266), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n239) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_U7 ( .A(
        Red_StateRegOutput[76]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n223), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n266) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_U6 ( .A(
        F_SD2_RedSB_inst_n59), .B(F_SD2_RedSB_inst_n60), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n223) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_U5 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n251), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n267) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_U4 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n222), .B(
        Red_StateRegOutput[74]), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n251) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_U3 ( .A(
        F_SD2_RedSB_inst_n59), .B(F_SD2_RedSB_inst_n58), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_76_n222) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_U69 ( .A(
        Red_StateRegOutput[78]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n280), .Z(Red_Feedback[35])
         );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_U68 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n279), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n278), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n280) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_U67 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n277), .B2(
        Red_StateRegOutput[79]), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n276), .C2(
        Red_StateRegOutput[82]), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n275), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n278) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_U66 ( .A1(
        Red_StateRegOutput[79]), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n277), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n276), .B2(
        Red_StateRegOutput[82]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n275) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_U65 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n274), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n273), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n276) );
  AOI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_U64 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n272), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n271), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n270), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n269), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n273) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_U63 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n268), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n267), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n266), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n265), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n264), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n269) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_U62 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n268), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n263), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n262), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n270) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_U61 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n268), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n263), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n261), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n262) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_U60 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n260), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n259), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n258), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n271) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_U59 ( .A(
        Red_StateRegOutput[77]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n257), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n274) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_U58 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n256), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n255), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n254), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n257) );
  OR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_U57 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n267), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n253), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n252), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n254) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_U56 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n251), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n250), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n249), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n252) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_U55 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n250), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n251), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n248), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n253) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_U54 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n247), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n246), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n245), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n244), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n255) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_U53 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n243), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n242), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n241), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n240), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n247) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_U52 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n239), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n238), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n240), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n237), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n236), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n277) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_U51 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n235), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n234), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n233), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n236) );
  AOI222_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_U50 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n251), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n249), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n251), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n232), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n249), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n232), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n234) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_U49 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n242), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n267), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n232) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_U48 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n263), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n246), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n249) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_U47 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n231), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n251) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_U46 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n256), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n230), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n237) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_U45 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n261), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n263), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n229), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n238) );
  NOR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_U44 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n267), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n244), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n259), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n229) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_U43 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n245), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n246), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n259) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_U42 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n268), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n228), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n244) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_U41 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n256), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n267) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_U40 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n242), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n245), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n261) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_U39 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n264), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n260), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n227), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n279) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_U38 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n246), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n226), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n225), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n227) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_U37 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n246), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n224), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n248), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n225) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_U36 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n235), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n248) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_U35 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n242), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n265), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n235) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_U34 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n239), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n228), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n265) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_U33 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n241), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n243), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n256), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n263), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n224) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_U32 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n240), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n245), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n243) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_U31 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n266), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n242), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n241) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_U30 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n272), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n223), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n258), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n226) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_U29 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n231), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n222), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n258) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_U28 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n240), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n228), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n223) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_U27 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n231), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n222), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n260) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_U26 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n228), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n256), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n222) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_U25 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n221), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n220), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n256) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_U24 ( .A(
        Red_StateRegOutput[77]), .B(F_SD2_RedSB_inst_n61), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n221) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_U23 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n263), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n228) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_U22 ( .A(
        Red_StateRegOutput[83]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n219), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n263) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_U21 ( .A(
        F_SD2_RedSB_inst_n64), .B(F_SD2_RedSB_inst_n63), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n219) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_U20 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n239), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n268), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n231) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_U19 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n266), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n268) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_U18 ( .A(
        Red_StateRegOutput[81]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n220), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n266) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_U17 ( .A(
        F_SD2_RedSB_inst_n62), .B(F_SD2_RedSB_inst_n63), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n220) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_U16 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n240), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n239) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_U15 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n218), .B(
        Red_StateRegOutput[80]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n240) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_U14 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n230), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n264) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_U13 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n250), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n246), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n230) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_U12 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n217), .B(
        F_SD2_RedSB_inst_n62), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n246) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_U11 ( .A(
        Red_StateRegOutput[78]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n218), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n217) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_U10 ( .A(
        F_SD2_RedSB_inst_n64), .B(F_SD2_RedSB_inst_n61), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n218) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_U9 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n242), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n245), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n250) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_U8 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n233), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n245) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_U7 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n216), .B(
        Red_StateRegOutput[79]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n233) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_U6 ( .A(
        F_SD2_RedSB_inst_n61), .B(F_SD2_RedSB_inst_n63), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n216) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_U5 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n272), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n242) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_U4 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n215), .B(
        F_SD2_RedSB_inst_n62), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n272) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_U3 ( .A(
        Red_StateRegOutput[82]), .B(F_SD2_RedSB_inst_n64), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_77_n215) );
  AOI222_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_U69 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n279), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n278), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n279), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n277), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n278), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n276), .ZN(Red_Feedback[36])
         );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_U68 ( .A(
        Red_StateRegOutput[82]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n275), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n276) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_U67 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n274), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n273), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n272), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n273), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n271), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n275) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_U66 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n270), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n269), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n268), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n269), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n267), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n271) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_U65 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n266), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n267) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_U64 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n265), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n264), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n268) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_U63 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n263), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n262), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n261), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n272) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_U62 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n260), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n259), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n262) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_U61 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n265), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n264), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n258), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n274) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_U60 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n265), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n264), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n257), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n258) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_U59 ( .A(
        Red_StateRegOutput[78]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n256), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n277) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_U58 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n255), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n254), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n253), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n256) );
  AOI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_U57 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n266), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n252), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n251), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n250), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n253) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_U56 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n249), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n248), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n260), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n261), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n250) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_U55 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n247), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n246), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n261) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_U54 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n245), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n260), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n244), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n243), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n249) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_U53 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n242), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n260) );
  NOR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_U52 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n241), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n240), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n239), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n251) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_U51 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n263), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n252) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_U50 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n247), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n246), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n263) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_U49 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n265), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n238), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n246) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_U48 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n244), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n238), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n254) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_U47 ( .A(
        Red_StateRegOutput[77]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n237), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n278) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_U46 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n238), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n236), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n235), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n237) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_U45 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n238), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n234), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n233), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n235) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_U44 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n244), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n247), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n259), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n248), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n233) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_U43 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n232), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n264), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n239), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n255), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n236) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_U42 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n257), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n241), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n255) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_U41 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n257), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n265), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n242), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n231), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n232) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_U40 ( .A(
        Red_StateRegOutput[79]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n230), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n279) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_U39 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n229), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n259), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n228), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n257), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n227), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n230) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_U38 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n226), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n225), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n224), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n223), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n227) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_U37 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n257), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n244), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n223) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_U36 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n222), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n224) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_U35 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n241), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n266), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n225) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_U34 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n257), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n239), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n266) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_U33 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n242), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n248), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n239) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_U32 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n259), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n257) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_U31 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n234), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n221), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n228) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_U30 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n222), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n247), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n231), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n240), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n221) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_U29 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n241), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n248), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n231) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_U28 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n273), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n248) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_U27 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n273), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n238), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n222) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_U26 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n273), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n245), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n244), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n247), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n234) );
  AND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_U25 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n270), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n264), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n247) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_U24 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n265), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n242), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n244) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_U23 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n240), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n265) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_U22 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n240), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n270), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n245) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_U21 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n241), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n270) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_U20 ( .A(
        Red_StateRegOutput[82]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n220), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n273) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_U19 ( .A(
        F_SD2_RedSB_inst_n63), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n219), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n259) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_U18 ( .A(
        Red_StateRegOutput[79]), .B(F_SD2_RedSB_inst_n61), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n219) );
  NOR4_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_U17 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n242), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n241), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n240), .A4(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n269), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n229) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_U16 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n243), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n269) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_U15 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n264), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n226), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n243) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_U14 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n238), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n226) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_U13 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n218), .B(
        Red_StateRegOutput[77]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n238) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_U12 ( .A(
        F_SD2_RedSB_inst_n61), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n217), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n218) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_U11 ( .A(
        Red_StateRegOutput[81]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n217), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n264) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_U10 ( .A(
        F_SD2_RedSB_inst_n63), .B(F_SD2_RedSB_inst_n62), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n217) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_U9 ( .A(
        Red_StateRegOutput[83]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n216), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n240) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_U8 ( .A(
        F_SD2_RedSB_inst_n63), .B(F_SD2_RedSB_inst_n64), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n216) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_U7 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n215), .B(
        Red_StateRegOutput[80]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n241) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_U6 ( .A(
        F_SD2_RedSB_inst_n61), .B(F_SD2_RedSB_inst_n64), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n215) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_U5 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n214), .B(
        Red_StateRegOutput[78]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n242) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_U4 ( .A(
        F_SD2_RedSB_inst_n61), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n220), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n214) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_U3 ( .A(
        F_SD2_RedSB_inst_n62), .B(F_SD2_RedSB_inst_n64), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_78_n220) );
  MUX2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_U54 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n240), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n239), .S(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n238), .Z(Red_Feedback[37])
         );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_U53 ( .A(
        Red_StateRegOutput[79]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n237), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n238) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_U52 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n236), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n235), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n234), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n233), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n237) );
  OR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_U51 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n232), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n231), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n230), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n233) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_U50 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n229), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n228), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n227), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n234) );
  AOI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_U49 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n226), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n225), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n224), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n223), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n236) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_U48 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n222), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n221), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n220), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n221), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n219), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n223) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_U47 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n226), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n225), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n218), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n221) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_U46 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n217), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n216), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n225) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_U45 ( .A(
        Red_StateRegOutput[82]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n215), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n239) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_U44 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n214), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n230), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n213), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n212), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n215) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_U43 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n228), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n226), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n211), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n232), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n212) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_U42 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n210), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n228), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n210), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n226), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n216), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n213) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_U41 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n220), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n216) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_U40 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n209), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n226) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_U39 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n208), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n207), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n228) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_U38 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n219), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n206), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n205), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n210) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_U37 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n219), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n206), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n208), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n205) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_U36 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n235), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n208) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_U35 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n222), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n204), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n229), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n214) );
  AND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_U34 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n206), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n219), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n204) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_U33 ( .A(
        Red_StateRegOutput[78]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n203), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n240) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_U32 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n202), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n201), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n200), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n201), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n199), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n203) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_U31 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n198), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n197), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n230), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n209), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n199) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_U30 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n227), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n220), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n218), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n197) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_U29 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n207), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n218) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_U28 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n222), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n201), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n227) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_U27 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n198), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n230), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n209), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n230), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n217), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n200) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_U26 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n231), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n206), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n209) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_U25 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n207), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n235), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n220), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n230) );
  AOI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_U24 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n229), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n211), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n207), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n224), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n198) );
  NOR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_U23 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n231), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n220), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n201), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n224) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_U22 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n219), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n220), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n211) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_U21 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n196), .B(
        Red_StateRegOutput[82]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n220) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_U20 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n201), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n219) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_U19 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n232), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n206), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n229) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_U18 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n195), .B(
        Red_StateRegOutput[81]), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n206) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_U17 ( .A(
        F_SD2_RedSB_inst_n63), .B(F_SD2_RedSB_inst_n62), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n195) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_U16 ( .A(
        Red_StateRegOutput[83]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n194), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n201) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_U15 ( .A(
        F_SD2_RedSB_inst_n63), .B(F_SD2_RedSB_inst_n64), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n194) );
  NOR4_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_U14 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n207), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n231), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n232), .A4(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n235), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n202) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_U13 ( .A(
        Red_StateRegOutput[79]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n193), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n235) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_U12 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n217), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n232) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_U11 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n192), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n193), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n217) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_U10 ( .A(
        F_SD2_RedSB_inst_n61), .B(F_SD2_RedSB_inst_n63), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n193) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_U9 ( .A(
        F_SD2_RedSB_inst_n62), .B(Red_StateRegOutput[77]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n192) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_U8 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n222), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n231) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_U7 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n191), .B(
        Red_StateRegOutput[80]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n222) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_U6 ( .A(
        F_SD2_RedSB_inst_n61), .B(F_SD2_RedSB_inst_n64), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n191) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_U5 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n190), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n196), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n207) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_U4 ( .A(
        F_SD2_RedSB_inst_n62), .B(F_SD2_RedSB_inst_n64), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n196) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_U3 ( .A(
        F_SD2_RedSB_inst_n61), .B(Red_StateRegOutput[78]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_79_n190) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_U71 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n289), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n291), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n290), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n288) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_U70 ( .A(
        Red_StateRegOutput[82]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n275), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n289) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_U69 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n274), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n273), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n272), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n276), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n275) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_U68 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n271), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n281), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n270), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n269), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n268), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n272) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_U67 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n267), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n266), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n285), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n265), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n270) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_U66 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n269), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n281) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_U65 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n280), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n279), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n271) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_U64 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n264), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n273) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_U63 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n263), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n262), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n261), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n274) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_U62 ( .A(
        Red_StateRegOutput[79]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n260), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n290) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_U61 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n259), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n269), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n258), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n257), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n260) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_U60 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n285), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n264), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n256), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n257) );
  NAND4_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_U59 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n261), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n255), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n283), .A4(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n269), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n258) );
  AOI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_U58 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n278), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n254), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n253), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n284), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n259) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_U57 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n265), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n266), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n252), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n284) );
  NOR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_U56 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n285), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n251), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n287), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n253) );
  AND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_U55 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n265), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n266), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n287) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_U54 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n250), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n266) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_U53 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n256), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n276), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n278) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_U52 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n252), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n267), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n247), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n248) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_U51 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n250), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n246), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n264), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n247) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_U50 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n283), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n286), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n264) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_U49 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n269), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n276), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n286) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_U48 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n251), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n263), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n252) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_U47 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n245), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n254), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n263) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_U46 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n244), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n249) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_U45 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n276), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n255), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n268), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n244) );
  AND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_U44 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n250), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n246), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n268) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_U43 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n285), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n279), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n246) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_U42 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n256), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n280), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n250) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_U41 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n262), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n280) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_U40 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n256), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n254), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n255) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_U39 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n282), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n262), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n261) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_U38 ( .A(
        Red_StateRegOutput[81]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n243), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n262) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_U37 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n285), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n282) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_U36 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n276), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n251) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_U35 ( .A(
        Red_StateRegOutput[82]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n242), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n276) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_U34 ( .A(
        F_SD2_RedSB_inst_n62), .B(F_SD2_RedSB_inst_n64), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n242) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_U33 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n269), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n245), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n277) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_U32 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n256), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n245) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_U31 ( .A(
        Red_StateRegOutput[80]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n241), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n256) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_U30 ( .A(
        F_SD2_RedSB_inst_n61), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n240), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n269) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_U29 ( .A(
        Red_StateRegOutput[79]), .B(F_SD2_RedSB_inst_n63), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n240) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_U28 ( .A(
        F_SD2_RedSB_inst_n62), .B(F_SD2_RedSB_inst_n63), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n243) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_U27 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n283), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n254), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n265) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_U26 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n279), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n254) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_U25 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n239), .B(
        Red_StateRegOutput[83]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n279) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_U24 ( .A(
        F_SD2_RedSB_inst_n63), .B(F_SD2_RedSB_inst_n64), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n239) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_U23 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n267), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n283) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_U22 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n238), .B(
        Red_StateRegOutput[78]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n267) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_U21 ( .A(
        F_SD2_RedSB_inst_n62), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n241), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n238) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_U20 ( .A(
        F_SD2_RedSB_inst_n61), .B(F_SD2_RedSB_inst_n64), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n241) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_U19 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n235), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n234), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n236), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n237), .ZN(Red_Feedback[38])
         );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_U18 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n235), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n230), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n234), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n237) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_U17 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n289), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n290), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n291), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n236) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_U16 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n289), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n290), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n288), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n235) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_U15 ( .A(
        Red_StateRegOutput[78]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n233), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n234) );
  AOI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_U14 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n267), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n249), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n232), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n248), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n233) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_U13 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n265), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n231), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n232) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_U12 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n261), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n251), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n277), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n285), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n231) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_U11 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n291), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n230) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_U10 ( .A(
        Red_StateRegOutput[77]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n229), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n285) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_U9 ( .A(
        F_SD2_RedSB_inst_n61), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n243), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n229) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_U8 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n228), .B(
        Red_StateRegOutput[77]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n291) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_U7 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n224), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n284), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n227), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n228) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_U6 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n283), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n225), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n282), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n226), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n227) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_U5 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n281), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n279), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n280), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n226) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_U4 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n276), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n277), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n280), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n278), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n225) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_U3 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n287), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n286), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n285), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_80_n224) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_U73 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n277), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n276), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n279), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n278) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_U72 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n275), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n274), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n273), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n277) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_U71 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n272), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n279) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_U70 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n267), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n266), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n265), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n268) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_U69 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n263), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n262), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n280) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_U68 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n265), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n281), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n261), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n276) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_U67 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n265), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n260), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n283) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_U66 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n263), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n264), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n258), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n285), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n259) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_U65 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n272), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n257), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n285) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_U64 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n270), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n256), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n282) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_U63 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n286), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n274) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_U62 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n260), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n255), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n286) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_U61 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n262), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n271), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n254), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n252) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_U60 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n273), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n251), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n250), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n253) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_U59 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n284), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n250) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_U58 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n270), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n256), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n284) );
  OR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_U57 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n275), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n257), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n256) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_U56 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n267), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n270) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_U55 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n258), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n275), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n251) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_U54 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n281), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n258) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_U53 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n272), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n248), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n247), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n249) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_U52 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n262), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n264), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n246), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n245), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n247) );
  OR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_U51 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n254), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n271), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n269), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n245) );
  OR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_U50 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n281), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n257), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n263), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n269) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_U49 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n260), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n254) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_U48 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n267), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n255), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n266), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n244), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n257), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n246) );
  AND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_U47 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n267), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n255), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n244) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_U46 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n275), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n260), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n266) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_U45 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n265), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n281), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n255) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_U44 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n263), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n265) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_U43 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n272), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n273), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n267) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_U42 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n273), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n257), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n264) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_U41 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n271), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n273) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_U40 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n275), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n281), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n262) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_U39 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n261), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n275) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_U38 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n261), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n243), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n263), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n243), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n257), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n248) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_U37 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n242), .B(
        Red_StateRegOutput[77]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n257) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_U36 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n241), .B(
        F_SD2_RedSB_inst_n62), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n242) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_U35 ( .A(
        Red_StateRegOutput[79]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n241), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n263) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_U34 ( .A(
        F_SD2_RedSB_inst_n63), .B(F_SD2_RedSB_inst_n61), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n241) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_U33 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n260), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n281), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n271), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n243) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_U32 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n240), .B(
        Red_StateRegOutput[80]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n271) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_U31 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n239), .B(
        F_SD2_RedSB_inst_n62), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n281) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_U30 ( .A(
        Red_StateRegOutput[82]), .B(F_SD2_RedSB_inst_n64), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n239) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_U29 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n238), .B(
        Red_StateRegOutput[78]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n260) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_U28 ( .A(
        F_SD2_RedSB_inst_n62), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n240), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n238) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_U27 ( .A(
        F_SD2_RedSB_inst_n61), .B(F_SD2_RedSB_inst_n64), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n240) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_U26 ( .A(
        Red_StateRegOutput[83]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n237), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n261) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_U25 ( .A(
        F_SD2_RedSB_inst_n63), .B(F_SD2_RedSB_inst_n64), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n237) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_U24 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n236), .B(
        Red_StateRegOutput[81]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n272) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_U23 ( .A(
        F_SD2_RedSB_inst_n63), .B(F_SD2_RedSB_inst_n62), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n236) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_U22 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n217), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n221), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n234), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n225), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n235), .ZN(Red_Feedback[39])
         );
  NOR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_U21 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n221), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n225), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n234), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n235) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_U20 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n232), .B2(
        Red_StateRegOutput[79]), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n233), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n234) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_U19 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n232), .B2(
        Red_StateRegOutput[79]), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n217), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n233) );
  AOI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_U18 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n271), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n227), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n229), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n231), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n232) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_U17 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n271), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n230), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n264), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n286), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n231) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_U16 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n280), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n230) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_U15 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n270), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n228), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n268), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n269), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n229) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_U14 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n266), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n228) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_U13 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n285), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n226), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n276), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n227) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_U12 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n275), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n283), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n226) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_U11 ( .A(
        Red_StateRegOutput[82]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n224), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n225) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_U10 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n285), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n286), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n222), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n223), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n224) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_U9 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n279), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n280), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n278), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n223) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_U8 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n284), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n282), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n284), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n283), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n281), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n222) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_U7 ( .A(
        Red_StateRegOutput[78]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n220), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n221) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_U6 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n219), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n218), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n220) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_U5 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n254), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n253), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n252), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n219) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_U4 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n266), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n259), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n282), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n274), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n218) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_U3 ( .A(
        Red_StateRegOutput[77]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n249), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_81_n217) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_U73 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n284), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n283), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n282), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n281), .ZN(Red_Feedback[40])
         );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_U72 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n280), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n281), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n279), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n283) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_U71 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n280), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n281), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n282), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n279) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_U70 ( .A(
        Red_StateRegOutput[82]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n278), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n282) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_U69 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n277), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n276), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n278) );
  NAND4_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_U68 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n275), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n274), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n273), .A4(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n272), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n276) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_U67 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n271), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n270), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n269), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n268), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n277) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_U66 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n267), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n268) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_U65 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n274), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n266), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n265), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n264), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n270) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_U64 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n263), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n265) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_U63 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n262), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n272), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n261), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n260), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n266) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_U62 ( .A(
        Red_StateRegOutput[78]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n259), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n281) );
  NOR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_U61 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n258), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n257), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n256), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n259) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_U60 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n255), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n254), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n255), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n253), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n252), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n256) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_U59 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n273), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n263), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n252) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_U58 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n251), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n250), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n263) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_U57 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n275), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n262), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n253) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_U56 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n271), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n269), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n254) );
  AOI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_U55 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n275), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n249), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n248), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n247), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n257) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_U54 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n246), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n245), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n275), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n247) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_U53 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n271), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n244), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n249) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_U52 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n245), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n271) );
  NOR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_U51 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n251), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n244), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n250), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n258) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_U50 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n260), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n248), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n250) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_U49 ( .A(
        Red_StateRegOutput[77]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n243), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n280) );
  AOI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_U48 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n275), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n242), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n241), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n240), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n243) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_U47 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n251), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n239), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n255), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n238), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n240) );
  OR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_U46 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n251), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n239), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n260), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n238) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_U45 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n237), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n248), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n244), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n255) );
  NOR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_U44 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n237), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n236), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n272), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n241) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_U43 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n274), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n262), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n246), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n235), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n236) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_U42 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n234), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n260), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n233), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n242) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_U41 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n232), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n246), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n262), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n233) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_U40 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n231), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n234) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_U39 ( .A(
        Red_StateRegOutput[79]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n230), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n284) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_U38 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n262), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n229), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n228), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n230) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_U37 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n267), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n227), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n226), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n264), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n228) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_U36 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n244), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n225), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n264) );
  NAND4_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_U35 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n237), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n269), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n274), .A4(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n227), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n226) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_U34 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n272), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n269) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_U33 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n237), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n273), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n262), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n231), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n267) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_U32 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n245), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n248), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n231) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_U31 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n244), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n239), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n273) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_U30 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n245), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n225), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n239) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_U29 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n260), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n237) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_U28 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n274), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n224), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n223), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n251), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n229) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_U27 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n232), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n244), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n261), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n244), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n235), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n224) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_U26 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n275), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n245), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n235) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_U25 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n227), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n275) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_U24 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n251), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n261) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_U23 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n227), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n272), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n251) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_U22 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n222), .B(
        Red_StateRegOutput[81]), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n272) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_U21 ( .A(
        F_SD2_RedSB_inst_n62), .B(F_SD2_RedSB_inst_n63), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n222) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_U20 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n221), .B(
        Red_StateRegOutput[80]), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n227) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_U19 ( .A(
        F_SD2_RedSB_inst_n61), .B(F_SD2_RedSB_inst_n64), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n221) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_U18 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n246), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n244) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_U17 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n220), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n219), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n246) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_U16 ( .A(
        F_SD2_RedSB_inst_n64), .B(Red_StateRegOutput[78]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n220) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_U15 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n223), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n232) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_U14 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n260), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n245), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n223) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_U13 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n218), .B(
        Red_StateRegOutput[82]), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n245) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_U12 ( .A(
        F_SD2_RedSB_inst_n62), .B(F_SD2_RedSB_inst_n64), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n218) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_U11 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n217), .B(
        F_SD2_RedSB_inst_n63), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n260) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_U10 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n219), .B(
        Red_StateRegOutput[77]), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n217) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_U9 ( .A(
        F_SD2_RedSB_inst_n61), .B(F_SD2_RedSB_inst_n62), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n219) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_U8 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n248), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n274) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_U7 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n216), .B(
        Red_StateRegOutput[83]), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n248) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_U6 ( .A(
        F_SD2_RedSB_inst_n63), .B(F_SD2_RedSB_inst_n64), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n216) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_U5 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n225), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n262) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_U4 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n215), .B(
        F_SD2_RedSB_inst_n63), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n225) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_U3 ( .A(
        Red_StateRegOutput[79]), .B(F_SD2_RedSB_inst_n61), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_82_n215) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_U65 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n283), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n282), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n281), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n280), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n279), .ZN(Red_Feedback[41])
         );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_U64 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n283), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n282), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n281), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n279) );
  MUX2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_U63 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n283), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n282), .S(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n278), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n280) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_U62 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n277), .B(
        Red_StateRegOutput[79]), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n278) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_U61 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n276), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n275), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n274), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n277) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_U60 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n273), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n274) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_U59 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n272), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n271), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n270), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n269), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n268), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n273) );
  AND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_U58 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n267), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n266), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n265), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n269) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_U57 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n266), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n264), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n263), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n262), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n275) );
  AOI222_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_U56 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n261), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n260), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n261), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n259), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n260), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n259), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n263) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_U55 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n258), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n268), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n259) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_U54 ( .A(
        Red_StateRegOutput[77]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n257), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n281) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_U53 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n268), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n256), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n255), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n257) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_U52 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n268), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n254), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n262), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n255) );
  AOI222_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_U51 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n261), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n260), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n261), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n253), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n260), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n253), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n254) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_U50 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n276), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n258), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n253) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_U49 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n252), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n251), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n250), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n249), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n256) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_U48 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n276), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n266), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n248), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n247), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n252) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_U47 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n264), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n247) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_U46 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n272), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n258), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n264) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_U45 ( .A(
        Red_StateRegOutput[78]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n246), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n282) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_U44 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n248), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n262), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n245), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n244), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n246) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_U43 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n248), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n243), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n244) );
  AOI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_U42 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n271), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n242), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n241), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n240), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n245) );
  NOR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_U41 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n270), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n239), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n250), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n240) );
  AND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_U40 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n238), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n268), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n260), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n241) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_U39 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n248), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n266), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n260) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_U38 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n251), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n237), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n249), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n238) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_U37 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n276), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n270), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n249) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_U36 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n258), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n236), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n262) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_U35 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n237), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n258) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_U34 ( .A(
        Red_StateRegOutput[82]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n235), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n283) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_U33 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n234), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n237), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n233), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n237), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n232), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n235) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_U32 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n251), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n268), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n267), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n236), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n271), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n232) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_U31 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n250), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n276), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n271) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_U30 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n237), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n248), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n250) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_U29 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n239), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n272), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n236) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_U28 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n242), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n265), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n243), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n233) );
  AND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_U27 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n261), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n231), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n243) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_U26 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n276), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n248), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n265) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_U25 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n230), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n229), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n248) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_U24 ( .A(
        F_SD2_RedSB_inst_n61), .B(Red_StateRegOutput[78]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n230) );
  OR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_U23 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n261), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n231), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n242) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_U22 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n268), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n266), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n231) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_U21 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n228), .B(
        Red_StateRegOutput[77]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n268) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_U20 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n227), .B(
        F_SD2_RedSB_inst_n62), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n228) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_U19 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n267), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n270), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n261) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_U18 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n272), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n270) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_U17 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n226), .B(
        Red_StateRegOutput[80]), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n272) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_U16 ( .A(
        F_SD2_RedSB_inst_n61), .B(F_SD2_RedSB_inst_n64), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n226) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_U15 ( .A(
        Red_StateRegOutput[82]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n229), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n237) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_U14 ( .A(
        F_SD2_RedSB_inst_n64), .B(F_SD2_RedSB_inst_n62), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n229) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_U13 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n225), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n234) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_U12 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n267), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n239), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n224), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n225) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_U11 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n267), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n239), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n276), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n224) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_U10 ( .A(
        Red_StateRegOutput[79]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n227), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n276) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_U9 ( .A(
        F_SD2_RedSB_inst_n63), .B(F_SD2_RedSB_inst_n61), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n227) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_U8 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n266), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n239) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_U7 ( .A(
        Red_StateRegOutput[83]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n223), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n266) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_U6 ( .A(
        F_SD2_RedSB_inst_n63), .B(F_SD2_RedSB_inst_n64), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n223) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_U5 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n251), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n267) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_U4 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n222), .B(
        Red_StateRegOutput[81]), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n251) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_U3 ( .A(
        F_SD2_RedSB_inst_n63), .B(F_SD2_RedSB_inst_n62), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_83_n222) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_U69 ( .A(
        Red_StateRegOutput[85]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n280), .Z(Red_Feedback[7]) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_U68 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n279), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n278), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n280) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_U67 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n277), .B2(
        Red_StateRegOutput[86]), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n276), .C2(
        Red_StateRegOutput[89]), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n275), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n278) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_U66 ( .A1(
        Red_StateRegOutput[86]), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n277), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n276), .B2(
        Red_StateRegOutput[89]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n275) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_U65 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n274), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n273), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n276) );
  AOI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_U64 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n272), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n271), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n270), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n269), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n273) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_U63 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n268), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n267), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n266), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n265), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n264), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n269) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_U62 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n268), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n263), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n262), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n270) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_U61 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n268), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n263), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n261), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n262) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_U60 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n260), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n259), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n258), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n271) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_U59 ( .A(
        Red_StateRegOutput[84]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n257), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n274) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_U58 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n253), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n252), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n251), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n254) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_U57 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n252), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n253), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n250), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n255) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_U56 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n242), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n241), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n243), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n240), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n239), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n277) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_U55 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n238), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n237), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n236), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n239) );
  AOI222_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_U54 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n253), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n251), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n253), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n235), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n251), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n235), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n237) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_U53 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n245), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n267), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n235) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_U52 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n263), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n249), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n251) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_U51 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n234), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n253) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_U50 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n256), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n233), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n240) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_U49 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n261), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n263), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n232), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n241) );
  NOR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_U48 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n267), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n247), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n259), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n232) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_U47 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n248), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n249), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n259) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_U46 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n268), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n231), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n247) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_U45 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n256), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n267) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_U44 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n245), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n248), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n261) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_U43 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n264), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n260), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n230), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n279) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_U42 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n249), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n229), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n228), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n230) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_U41 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n249), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n227), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n250), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n228) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_U40 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n238), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n250) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_U39 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n245), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n265), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n238) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_U38 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n242), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n231), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n265) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_U37 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n244), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n246), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n256), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n263), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n227) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_U36 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n243), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n248), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n246) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_U35 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n266), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n245), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n244) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_U34 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n272), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n226), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n258), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n229) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_U33 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n234), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n225), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n258) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_U32 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n243), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n231), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n226) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_U31 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n234), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n225), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n260) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_U30 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n231), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n256), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n225) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_U29 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n224), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n223), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n256) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_U28 ( .A(
        Red_StateRegOutput[84]), .B(F_SD2_RedSB_inst_n65), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n224) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_U27 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n263), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n231) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_U26 ( .A(
        Red_StateRegOutput[90]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n222), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n263) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_U25 ( .A(
        F_SD2_RedSB_inst_n68), .B(F_SD2_RedSB_inst_n67), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n222) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_U24 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n242), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n268), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n234) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_U23 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n266), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n268) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_U22 ( .A(
        Red_StateRegOutput[88]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n223), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n266) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_U21 ( .A(
        F_SD2_RedSB_inst_n66), .B(F_SD2_RedSB_inst_n67), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n223) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_U20 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n243), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n242) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_U19 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n221), .B(
        Red_StateRegOutput[87]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n243) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_U18 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n233), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n264) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_U17 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n252), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n249), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n233) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_U16 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n220), .B(
        F_SD2_RedSB_inst_n66), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n249) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_U15 ( .A(
        Red_StateRegOutput[85]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n221), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n220) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_U14 ( .A(
        F_SD2_RedSB_inst_n68), .B(F_SD2_RedSB_inst_n65), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n221) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_U13 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n245), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n248), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n252) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_U12 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n236), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n248) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_U11 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n219), .B(
        Red_StateRegOutput[86]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n236) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_U10 ( .A(
        F_SD2_RedSB_inst_n65), .B(F_SD2_RedSB_inst_n67), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n219) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_U9 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n272), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n245) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_U8 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n218), .B(
        F_SD2_RedSB_inst_n66), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n272) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_U7 ( .A(
        Red_StateRegOutput[89]), .B(F_SD2_RedSB_inst_n68), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n218) );
  OAI33_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_U6 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n256), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n215), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n217), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n267), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n255), .B3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n254), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n257) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_U5 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n249), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n216), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n217) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_U4 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n245), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n246), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n243), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n244), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n216) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_U3 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n248), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n247), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_84_n215) );
  AOI222_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_U69 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n279), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n278), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n279), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n277), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n278), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n276), .ZN(Red_Feedback[8])
         );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_U68 ( .A(
        Red_StateRegOutput[89]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n275), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n276) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_U67 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n274), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n273), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n272), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n273), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n271), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n275) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_U66 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n270), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n269), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n268), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n269), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n267), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n271) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_U65 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n266), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n267) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_U64 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n265), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n264), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n268) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_U63 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n263), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n262), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n261), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n272) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_U62 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n260), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n259), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n262) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_U61 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n265), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n264), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n258), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n274) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_U60 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n265), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n264), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n257), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n258) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_U59 ( .A(
        Red_StateRegOutput[85]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n256), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n277) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_U58 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n255), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n254), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n253), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n256) );
  AOI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_U57 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n266), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n252), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n251), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n250), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n253) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_U56 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n249), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n248), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n260), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n261), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n250) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_U55 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n247), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n246), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n261) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_U54 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n245), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n260), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n244), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n243), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n249) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_U53 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n242), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n260) );
  NOR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_U52 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n241), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n240), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n239), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n251) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_U51 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n263), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n252) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_U50 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n247), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n246), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n263) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_U49 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n265), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n238), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n246) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_U48 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n244), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n238), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n254) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_U47 ( .A(
        Red_StateRegOutput[84]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n237), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n278) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_U46 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n238), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n236), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n235), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n237) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_U45 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n238), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n234), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n233), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n235) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_U44 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n244), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n247), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n259), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n248), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n233) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_U43 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n232), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n264), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n239), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n255), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n236) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_U42 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n257), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n241), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n255) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_U41 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n257), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n265), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n242), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n231), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n232) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_U40 ( .A(
        Red_StateRegOutput[86]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n230), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n279) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_U39 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n229), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n259), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n228), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n257), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n227), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n230) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_U38 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n226), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n225), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n224), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n223), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n227) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_U37 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n257), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n244), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n223) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_U36 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n222), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n224) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_U35 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n241), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n266), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n225) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_U34 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n257), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n239), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n266) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_U33 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n242), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n248), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n239) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_U32 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n259), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n257) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_U31 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n234), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n221), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n228) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_U30 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n222), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n247), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n231), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n240), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n221) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_U29 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n241), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n248), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n231) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_U28 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n273), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n248) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_U27 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n273), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n238), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n222) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_U26 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n273), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n245), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n244), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n247), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n234) );
  AND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_U25 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n270), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n264), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n247) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_U24 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n265), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n242), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n244) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_U23 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n240), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n265) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_U22 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n240), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n270), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n245) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_U21 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n241), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n270) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_U20 ( .A(
        Red_StateRegOutput[89]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n220), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n273) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_U19 ( .A(
        F_SD2_RedSB_inst_n67), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n219), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n259) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_U18 ( .A(
        Red_StateRegOutput[86]), .B(F_SD2_RedSB_inst_n65), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n219) );
  NOR4_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_U17 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n242), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n241), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n240), .A4(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n269), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n229) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_U16 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n243), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n269) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_U15 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n264), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n226), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n243) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_U14 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n238), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n226) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_U13 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n218), .B(
        Red_StateRegOutput[84]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n238) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_U12 ( .A(
        F_SD2_RedSB_inst_n65), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n217), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n218) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_U11 ( .A(
        Red_StateRegOutput[88]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n217), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n264) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_U10 ( .A(
        F_SD2_RedSB_inst_n67), .B(F_SD2_RedSB_inst_n66), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n217) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_U9 ( .A(
        Red_StateRegOutput[90]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n216), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n240) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_U8 ( .A(
        F_SD2_RedSB_inst_n67), .B(F_SD2_RedSB_inst_n68), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n216) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_U7 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n215), .B(
        Red_StateRegOutput[87]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n241) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_U6 ( .A(
        F_SD2_RedSB_inst_n65), .B(F_SD2_RedSB_inst_n68), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n215) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_U5 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n214), .B(
        Red_StateRegOutput[85]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n242) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_U4 ( .A(
        F_SD2_RedSB_inst_n65), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n220), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n214) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_U3 ( .A(
        F_SD2_RedSB_inst_n66), .B(F_SD2_RedSB_inst_n68), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_85_n220) );
  MUX2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_U54 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n240), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n239), .S(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n238), .Z(Red_Feedback[9]) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_U53 ( .A(
        Red_StateRegOutput[86]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n237), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n238) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_U52 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n236), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n235), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n234), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n233), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n237) );
  OR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_U51 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n232), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n231), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n230), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n233) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_U50 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n229), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n228), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n227), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n234) );
  AOI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_U49 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n226), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n225), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n224), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n223), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n236) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_U48 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n222), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n221), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n220), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n221), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n219), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n223) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_U47 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n226), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n225), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n218), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n221) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_U46 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n217), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n216), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n225) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_U45 ( .A(
        Red_StateRegOutput[89]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n215), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n239) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_U44 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n214), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n230), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n213), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n212), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n215) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_U43 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n228), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n226), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n211), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n232), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n212) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_U42 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n210), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n228), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n210), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n226), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n216), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n213) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_U41 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n220), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n216) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_U40 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n209), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n226) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_U39 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n208), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n207), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n228) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_U38 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n219), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n206), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n205), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n210) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_U37 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n219), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n206), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n208), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n205) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_U36 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n235), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n208) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_U35 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n222), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n204), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n229), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n214) );
  AND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_U34 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n206), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n219), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n204) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_U33 ( .A(
        Red_StateRegOutput[85]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n203), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n240) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_U32 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n202), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n201), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n200), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n201), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n199), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n203) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_U31 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n198), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n197), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n230), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n209), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n199) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_U30 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n227), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n220), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n218), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n197) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_U29 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n207), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n218) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_U28 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n222), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n201), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n227) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_U27 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n198), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n230), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n209), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n230), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n217), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n200) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_U26 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n231), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n206), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n209) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_U25 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n207), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n235), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n220), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n230) );
  AOI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_U24 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n229), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n211), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n207), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n224), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n198) );
  NOR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_U23 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n231), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n220), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n201), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n224) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_U22 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n219), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n220), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n211) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_U21 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n196), .B(
        Red_StateRegOutput[89]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n220) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_U20 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n201), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n219) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_U19 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n232), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n206), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n229) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_U18 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n195), .B(
        Red_StateRegOutput[88]), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n206) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_U17 ( .A(
        F_SD2_RedSB_inst_n67), .B(F_SD2_RedSB_inst_n66), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n195) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_U16 ( .A(
        Red_StateRegOutput[90]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n194), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n201) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_U15 ( .A(
        F_SD2_RedSB_inst_n67), .B(F_SD2_RedSB_inst_n68), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n194) );
  NOR4_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_U14 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n207), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n231), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n232), .A4(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n235), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n202) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_U13 ( .A(
        Red_StateRegOutput[86]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n193), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n235) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_U12 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n217), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n232) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_U11 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n192), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n193), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n217) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_U10 ( .A(
        F_SD2_RedSB_inst_n65), .B(F_SD2_RedSB_inst_n67), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n193) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_U9 ( .A(
        F_SD2_RedSB_inst_n66), .B(Red_StateRegOutput[84]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n192) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_U8 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n222), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n231) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_U7 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n191), .B(
        Red_StateRegOutput[87]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n222) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_U6 ( .A(
        F_SD2_RedSB_inst_n65), .B(F_SD2_RedSB_inst_n68), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n191) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_U5 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n190), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n196), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n207) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_U4 ( .A(
        F_SD2_RedSB_inst_n66), .B(F_SD2_RedSB_inst_n68), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n196) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_U3 ( .A(
        F_SD2_RedSB_inst_n65), .B(Red_StateRegOutput[85]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_86_n190) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_U70 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n290), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n289), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n288), .ZN(Red_Feedback[10])
         );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_U69 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n290), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n287), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n288) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_U68 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n286), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n285), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n284), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n287) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_U67 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n283), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n282), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n286), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n284) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_U66 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n289), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n285) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_U65 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n283), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n282), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n281), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n289) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_U64 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n282), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n286), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n283), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n281) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_U63 ( .A(
        Red_StateRegOutput[89]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n268), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n282) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_U62 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n267), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n266), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n265), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n269), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n268) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_U61 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n264), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n274), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n263), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n262), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n261), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n265) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_U60 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n260), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n259), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n278), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n258), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n263) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_U59 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n262), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n274) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_U58 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n273), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n272), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n264) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_U57 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n257), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n266) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_U56 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n256), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n255), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n254), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n267) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_U55 ( .A(
        Red_StateRegOutput[86]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n253), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n283) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_U54 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n252), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n262), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n251), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n250), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n253) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_U53 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n278), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n257), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n249), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n250) );
  NAND4_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_U52 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n254), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n248), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n276), .A4(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n262), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n251) );
  AOI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_U51 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n271), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n247), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n246), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n277), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n252) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_U50 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n258), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n259), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n245), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n277) );
  NOR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_U49 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n278), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n244), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n280), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n246) );
  AND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_U48 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n258), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n259), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n280) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_U47 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n243), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n259) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_U46 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n249), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n269), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n271) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_U45 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n242), .B(
        Red_StateRegOutput[85]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n290) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_U44 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n276), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n279), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n257) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_U43 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n262), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n269), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n279) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_U42 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n244), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n256), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n245) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_U41 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n240), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n247), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n256) );
  AND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_U40 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n243), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n241), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n261) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_U39 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n278), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n272), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n241) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_U38 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n249), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n273), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n243) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_U37 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n255), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n273) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_U36 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n249), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n247), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n248) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_U35 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n275), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n255), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n254) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_U34 ( .A(
        Red_StateRegOutput[88]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n239), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n255) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_U33 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n278), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n275) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_U32 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n269), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n244) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_U31 ( .A(
        Red_StateRegOutput[89]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n238), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n269) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_U30 ( .A(
        F_SD2_RedSB_inst_n66), .B(F_SD2_RedSB_inst_n68), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n238) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_U29 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n262), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n240), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n270) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_U28 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n249), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n240) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_U27 ( .A(
        Red_StateRegOutput[87]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n237), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n249) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_U26 ( .A(
        F_SD2_RedSB_inst_n65), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n236), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n262) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_U25 ( .A(
        Red_StateRegOutput[86]), .B(F_SD2_RedSB_inst_n67), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n236) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_U24 ( .A(
        F_SD2_RedSB_inst_n66), .B(F_SD2_RedSB_inst_n67), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n239) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_U23 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n276), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n247), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n258) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_U22 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n272), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n247) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_U21 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n235), .B(
        Red_StateRegOutput[90]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n272) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_U20 ( .A(
        F_SD2_RedSB_inst_n67), .B(F_SD2_RedSB_inst_n68), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n235) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_U19 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n260), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n276) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_U18 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n234), .B(
        Red_StateRegOutput[85]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n260) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_U17 ( .A(
        F_SD2_RedSB_inst_n66), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n237), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n234) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_U16 ( .A(
        F_SD2_RedSB_inst_n65), .B(F_SD2_RedSB_inst_n68), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n237) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_U15 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n258), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n230), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n232), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n233), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n242) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_U14 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n261), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n269), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n261), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n248), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n260), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n233) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_U13 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n243), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n257), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n241), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n257), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n231), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n232) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_U12 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n260), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n245), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n231) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_U11 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n278), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n270), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n244), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n254), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n230) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_U10 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n229), .B(
        Red_StateRegOutput[84]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n286) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_U9 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n225), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n277), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n228), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n229) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_U8 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n276), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n226), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n275), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n227), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n228) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_U7 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n274), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n272), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n273), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n227) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_U6 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n269), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n270), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n273), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n271), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n226) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_U5 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n280), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n279), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n278), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n225) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_U4 ( .A(
        Red_StateRegOutput[84]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n224), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n278) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_U3 ( .A(
        F_SD2_RedSB_inst_n65), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n239), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_87_n224) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_U73 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n282), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n281), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n282), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n280), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n279), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n283) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_U72 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n278), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n277), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n276), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n284) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_U71 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n275), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n274), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n277), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n276) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_U70 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n273), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n272), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n271), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n275) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_U69 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n270), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n277) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_U68 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n264), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n263), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n262), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n265) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_U67 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n263), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n267) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_U66 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n278), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n261) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_U65 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n259), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n258), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n278) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_U64 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n262), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n279), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n256), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n274) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_U63 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n281), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n273), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n257) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_U62 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n262), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n255), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n281) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_U61 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n272), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n280), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n263), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n252), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n253) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_U60 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n259), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n260), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n251), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n285), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n252) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_U59 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n270), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n250), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n285) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_U58 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n268), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n249), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n280) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_U57 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n286), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n272) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_U56 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n255), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n248), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n286) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_U55 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n247), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n246), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n245), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n254) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_U54 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n258), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n269), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n247), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n245) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_U53 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n271), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n244), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n243), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n246) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_U52 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n282), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n243) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_U51 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n268), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n249), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n282) );
  OR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_U50 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n273), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n250), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n249) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_U49 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n264), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n268) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_U48 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n251), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n273), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n244) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_U47 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n279), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n251) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_U46 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n270), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n241), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n240), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n242) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_U45 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n258), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n260), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n239), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n238), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n240) );
  OR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_U44 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n247), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n269), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n266), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n238) );
  OR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_U43 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n279), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n250), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n259), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n266) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_U42 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n255), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n247) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_U41 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n264), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n248), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n263), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n237), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n250), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n239) );
  AND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_U40 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n264), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n248), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n237) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_U39 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n273), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n255), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n263) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_U38 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n262), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n279), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n248) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_U37 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n259), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n262) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_U36 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n270), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n271), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n264) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_U35 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n271), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n250), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n260) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_U34 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n269), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n271) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_U33 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n273), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n279), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n258) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_U32 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n256), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n273) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_U31 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n256), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n236), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n259), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n236), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n250), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n241) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_U30 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n235), .B(
        Red_StateRegOutput[84]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n250) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_U29 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n234), .B(
        F_SD2_RedSB_inst_n66), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n235) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_U28 ( .A(
        Red_StateRegOutput[86]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n234), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n259) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_U27 ( .A(
        F_SD2_RedSB_inst_n67), .B(F_SD2_RedSB_inst_n65), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n234) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_U26 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n255), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n279), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n269), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n236) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_U25 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n233), .B(
        Red_StateRegOutput[87]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n269) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_U24 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n232), .B(
        F_SD2_RedSB_inst_n66), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n279) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_U23 ( .A(
        Red_StateRegOutput[89]), .B(F_SD2_RedSB_inst_n68), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n232) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_U22 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n231), .B(
        Red_StateRegOutput[85]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n255) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_U21 ( .A(
        F_SD2_RedSB_inst_n66), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n233), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n231) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_U20 ( .A(
        F_SD2_RedSB_inst_n65), .B(F_SD2_RedSB_inst_n68), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n233) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_U19 ( .A(
        Red_StateRegOutput[90]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n230), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n256) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_U18 ( .A(
        F_SD2_RedSB_inst_n67), .B(F_SD2_RedSB_inst_n68), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n230) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_U17 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n229), .B(
        Red_StateRegOutput[88]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n270) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_U16 ( .A(
        F_SD2_RedSB_inst_n67), .B(F_SD2_RedSB_inst_n66), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n229) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_U15 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n217), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n219), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n227), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n221), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n228), .ZN(Red_Feedback[11])
         );
  NOR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_U14 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n219), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n221), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n227), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n228) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_U13 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n225), .B2(
        Red_StateRegOutput[86]), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n226), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n227) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_U12 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n225), .B2(
        Red_StateRegOutput[86]), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n217), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n226) );
  AOI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_U11 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n269), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n222), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n223), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n224), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n225) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_U10 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n286), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n260), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n261), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n269), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n224) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_U9 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n265), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n266), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n267), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n268), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n223) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_U8 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n285), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n257), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n274), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n222) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_U7 ( .A(
        Red_StateRegOutput[89]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n220), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n221) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_U6 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n286), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n285), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n284), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n283), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n220) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_U5 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n218), .B(
        Red_StateRegOutput[85]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n219) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_U4 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n254), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n253), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n218) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_U3 ( .A(
        Red_StateRegOutput[84]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n242), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_88_n217) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_U72 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n283), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n282), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n281), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n280), .ZN(Red_Feedback[12])
         );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_U71 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n279), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n280), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n278), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n282) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_U70 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n279), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n280), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n281), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n278) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_U69 ( .A(
        Red_StateRegOutput[89]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n277), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n281) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_U68 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n276), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n275), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n277) );
  NAND4_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_U67 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n274), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n273), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n272), .A4(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n271), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n275) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_U66 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n270), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n269), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n268), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n267), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n276) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_U65 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n266), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n267) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_U64 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n273), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n265), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n264), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n263), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n269) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_U63 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n262), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n264) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_U62 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n261), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n271), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n260), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n259), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n265) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_U61 ( .A(
        Red_StateRegOutput[85]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n258), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n280) );
  NOR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_U60 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n257), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n256), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n255), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n258) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_U59 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n253), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n252), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n262) );
  AOI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_U58 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n274), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n251), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n250), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n249), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n256) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_U57 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n248), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n247), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n274), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n249) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_U56 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n270), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n246), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n251) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_U55 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n247), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n270) );
  NOR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_U54 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n253), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n246), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n252), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n257) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_U53 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n259), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n250), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n252) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_U52 ( .A(
        Red_StateRegOutput[84]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n245), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n279) );
  AOI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_U51 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n274), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n244), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n243), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n242), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n245) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_U50 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n253), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n241), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n254), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n240), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n242) );
  OR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_U49 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n253), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n241), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n259), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n240) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_U48 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n239), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n250), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n246), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n254) );
  NOR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_U47 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n239), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n238), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n271), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n243) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_U46 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n273), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n261), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n248), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n237), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n238) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_U45 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n236), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n259), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n235), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n244) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_U44 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n234), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n248), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n261), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n235) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_U43 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n233), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n236) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_U42 ( .A(
        Red_StateRegOutput[86]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n232), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n283) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_U41 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n261), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n231), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n230), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n232) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_U40 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n266), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n229), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n228), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n263), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n230) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_U39 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n246), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n227), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n263) );
  NAND4_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_U38 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n239), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n268), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n273), .A4(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n229), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n228) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_U37 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n271), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n268) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_U36 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n239), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n272), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n261), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n233), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n266) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_U35 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n247), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n250), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n233) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_U34 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n246), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n241), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n272) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_U33 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n247), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n227), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n241) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_U32 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n259), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n239) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_U31 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n273), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n226), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n225), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n253), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n231) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_U30 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n234), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n246), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n260), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n246), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n237), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n226) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_U29 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n274), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n247), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n237) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_U28 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n229), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n274) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_U27 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n253), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n260) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_U26 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n229), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n271), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n253) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_U25 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n224), .B(
        Red_StateRegOutput[88]), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n271) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_U24 ( .A(
        F_SD2_RedSB_inst_n66), .B(F_SD2_RedSB_inst_n67), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n224) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_U23 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n223), .B(
        Red_StateRegOutput[87]), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n229) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_U22 ( .A(
        F_SD2_RedSB_inst_n65), .B(F_SD2_RedSB_inst_n68), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n223) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_U21 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n248), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n246) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_U20 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n222), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n221), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n248) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_U19 ( .A(
        F_SD2_RedSB_inst_n68), .B(Red_StateRegOutput[85]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n222) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_U18 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n225), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n234) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_U17 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n259), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n247), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n225) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_U16 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n220), .B(
        Red_StateRegOutput[89]), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n247) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_U15 ( .A(
        F_SD2_RedSB_inst_n66), .B(F_SD2_RedSB_inst_n68), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n220) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_U14 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n219), .B(
        F_SD2_RedSB_inst_n67), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n259) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_U13 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n221), .B(
        Red_StateRegOutput[84]), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n219) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_U12 ( .A(
        F_SD2_RedSB_inst_n65), .B(F_SD2_RedSB_inst_n66), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n221) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_U11 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n250), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n273) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_U10 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n218), .B(
        Red_StateRegOutput[90]), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n250) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_U9 ( .A(
        F_SD2_RedSB_inst_n67), .B(F_SD2_RedSB_inst_n68), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n218) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_U8 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n227), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n261) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_U7 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n217), .B(
        F_SD2_RedSB_inst_n67), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n227) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_U6 ( .A(
        Red_StateRegOutput[86]), .B(F_SD2_RedSB_inst_n65), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n217) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_U5 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n254), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n215), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n216), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n255) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_U4 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n272), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n262), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n216) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_U3 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n268), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n270), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n261), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n274), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_89_n215) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_U65 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n283), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n282), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n281), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n280), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n279), .ZN(Red_Feedback[13])
         );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_U64 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n283), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n282), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n281), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n279) );
  MUX2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_U63 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n283), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n282), .S(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n278), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n280) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_U62 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n277), .B(
        Red_StateRegOutput[86]), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n278) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_U61 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n276), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n275), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n274), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n277) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_U60 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n273), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n274) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_U59 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n272), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n271), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n270), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n269), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n268), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n273) );
  AND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_U58 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n267), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n266), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n265), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n269) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_U57 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n266), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n264), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n263), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n262), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n275) );
  AOI222_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_U56 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n261), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n260), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n261), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n259), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n260), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n259), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n263) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_U55 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n258), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n268), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n259) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_U54 ( .A(
        Red_StateRegOutput[84]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n257), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n281) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_U53 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n268), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n256), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n255), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n257) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_U52 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n268), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n254), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n262), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n255) );
  AOI222_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_U51 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n261), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n260), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n261), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n253), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n260), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n253), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n254) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_U50 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n276), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n258), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n253) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_U49 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n252), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n251), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n250), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n249), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n256) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_U48 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n276), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n266), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n248), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n247), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n252) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_U47 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n264), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n247) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_U46 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n272), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n258), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n264) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_U45 ( .A(
        Red_StateRegOutput[85]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n246), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n282) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_U44 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n248), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n262), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n245), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n244), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n246) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_U43 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n248), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n243), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n244) );
  AOI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_U42 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n271), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n242), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n241), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n240), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n245) );
  NOR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_U41 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n270), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n239), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n250), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n240) );
  AND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_U40 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n238), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n268), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n260), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n241) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_U39 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n248), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n266), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n260) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_U38 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n251), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n237), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n249), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n238) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_U37 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n276), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n270), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n249) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_U36 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n258), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n236), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n262) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_U35 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n237), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n258) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_U34 ( .A(
        Red_StateRegOutput[89]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n235), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n283) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_U33 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n234), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n237), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n233), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n237), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n232), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n235) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_U32 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n251), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n268), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n267), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n236), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n271), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n232) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_U31 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n250), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n276), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n271) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_U30 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n237), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n248), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n250) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_U29 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n239), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n272), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n236) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_U28 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n242), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n265), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n243), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n233) );
  AND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_U27 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n261), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n231), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n243) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_U26 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n276), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n248), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n265) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_U25 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n230), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n229), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n248) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_U24 ( .A(
        F_SD2_RedSB_inst_n65), .B(Red_StateRegOutput[85]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n230) );
  OR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_U23 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n261), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n231), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n242) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_U22 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n268), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n266), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n231) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_U21 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n228), .B(
        Red_StateRegOutput[84]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n268) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_U20 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n227), .B(
        F_SD2_RedSB_inst_n66), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n228) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_U19 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n267), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n270), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n261) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_U18 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n272), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n270) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_U17 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n226), .B(
        Red_StateRegOutput[87]), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n272) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_U16 ( .A(
        F_SD2_RedSB_inst_n65), .B(F_SD2_RedSB_inst_n68), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n226) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_U15 ( .A(
        Red_StateRegOutput[89]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n229), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n237) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_U14 ( .A(
        F_SD2_RedSB_inst_n68), .B(F_SD2_RedSB_inst_n66), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n229) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_U13 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n225), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n234) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_U12 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n267), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n239), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n224), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n225) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_U11 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n267), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n239), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n276), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n224) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_U10 ( .A(
        Red_StateRegOutput[86]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n227), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n276) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_U9 ( .A(
        F_SD2_RedSB_inst_n67), .B(F_SD2_RedSB_inst_n65), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n227) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_U8 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n266), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n239) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_U7 ( .A(
        Red_StateRegOutput[90]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n223), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n266) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_U6 ( .A(
        F_SD2_RedSB_inst_n67), .B(F_SD2_RedSB_inst_n68), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n223) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_U5 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n251), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n267) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_U4 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n222), .B(
        Red_StateRegOutput[88]), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n251) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_U3 ( .A(
        F_SD2_RedSB_inst_n67), .B(F_SD2_RedSB_inst_n66), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_90_n222) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_U69 ( .A(
        Red_StateRegOutput[92]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n280), .Z(Red_Feedback[14])
         );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_U68 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n279), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n278), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n280) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_U67 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n277), .B2(
        Red_StateRegOutput[93]), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n276), .C2(
        Red_StateRegOutput[96]), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n275), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n278) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_U66 ( .A1(
        Red_StateRegOutput[93]), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n277), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n276), .B2(
        Red_StateRegOutput[96]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n275) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_U65 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n274), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n273), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n276) );
  AOI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_U64 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n272), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n271), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n270), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n269), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n273) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_U63 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n268), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n267), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n266), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n265), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n264), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n269) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_U62 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n268), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n263), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n262), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n270) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_U61 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n268), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n263), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n261), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n262) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_U60 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n260), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n259), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n258), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n271) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_U59 ( .A(
        Red_StateRegOutput[91]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n257), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n274) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_U58 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n253), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n252), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n251), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n254) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_U57 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n252), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n253), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n250), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n255) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_U56 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n245), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n244), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n243), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n242), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n249) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_U55 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n241), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n240), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n242), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n239), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n238), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n277) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_U54 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n237), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n236), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n235), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n238) );
  AOI222_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_U53 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n253), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n251), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n253), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n234), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n251), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n234), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n236) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_U52 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n244), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n267), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n234) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_U51 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n263), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n248), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n251) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_U50 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n233), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n253) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_U49 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n256), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n232), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n239) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_U48 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n261), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n263), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n231), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n240) );
  NOR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_U47 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n267), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n246), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n259), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n231) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_U46 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n247), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n248), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n259) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_U45 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n268), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n230), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n246) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_U44 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n256), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n267) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_U43 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n244), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n247), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n261) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_U42 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n264), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n260), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n229), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n279) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_U41 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n248), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n228), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n227), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n229) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_U40 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n248), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n226), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n250), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n227) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_U39 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n237), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n250) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_U38 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n244), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n265), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n237) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_U37 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n241), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n230), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n265) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_U36 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n243), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n245), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n256), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n263), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n226) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_U35 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n242), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n247), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n245) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_U34 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n266), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n244), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n243) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_U33 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n272), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n225), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n258), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n228) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_U32 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n233), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n224), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n258) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_U31 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n242), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n230), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n225) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_U30 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n233), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n224), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n260) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_U29 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n230), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n256), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n224) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_U28 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n223), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n222), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n256) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_U27 ( .A(
        Red_StateRegOutput[91]), .B(F_SD2_RedSB_inst_n69), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n223) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_U26 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n263), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n230) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_U25 ( .A(
        Red_StateRegOutput[97]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n221), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n263) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_U24 ( .A(
        F_SD2_RedSB_inst_n72), .B(F_SD2_RedSB_inst_n71), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n221) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_U23 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n241), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n268), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n233) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_U22 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n266), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n268) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_U21 ( .A(
        Red_StateRegOutput[95]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n222), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n266) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_U20 ( .A(
        F_SD2_RedSB_inst_n70), .B(F_SD2_RedSB_inst_n71), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n222) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_U19 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n242), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n241) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_U18 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n220), .B(
        Red_StateRegOutput[94]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n242) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_U17 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n232), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n264) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_U16 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n252), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n248), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n232) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_U15 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n219), .B(
        F_SD2_RedSB_inst_n70), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n248) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_U14 ( .A(
        Red_StateRegOutput[92]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n220), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n219) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_U13 ( .A(
        F_SD2_RedSB_inst_n72), .B(F_SD2_RedSB_inst_n69), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n220) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_U12 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n244), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n247), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n252) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_U11 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n235), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n247) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_U10 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n218), .B(
        Red_StateRegOutput[93]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n235) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_U9 ( .A(
        F_SD2_RedSB_inst_n69), .B(F_SD2_RedSB_inst_n71), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n218) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_U8 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n272), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n244) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_U7 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n217), .B(
        F_SD2_RedSB_inst_n70), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n272) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_U6 ( .A(
        Red_StateRegOutput[96]), .B(F_SD2_RedSB_inst_n72), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n217) );
  OAI33_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_U5 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n256), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n215), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n216), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n267), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n255), .B3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n254), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n257) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_U4 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n249), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n248), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n216) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_U3 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n247), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n246), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_91_n215) );
  AOI222_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_U69 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n279), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n278), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n279), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n277), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n278), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n276), .ZN(Red_Feedback[15])
         );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_U68 ( .A(
        Red_StateRegOutput[96]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n275), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n276) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_U67 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n274), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n273), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n272), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n273), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n271), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n275) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_U66 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n270), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n269), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n268), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n269), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n267), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n271) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_U65 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n266), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n267) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_U64 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n265), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n264), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n268) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_U63 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n263), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n262), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n261), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n272) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_U62 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n260), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n259), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n262) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_U61 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n265), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n264), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n258), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n274) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_U60 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n265), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n264), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n257), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n258) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_U59 ( .A(
        Red_StateRegOutput[92]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n256), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n277) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_U58 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n255), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n254), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n253), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n256) );
  AOI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_U57 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n266), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n252), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n251), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n250), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n253) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_U56 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n249), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n248), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n260), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n261), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n250) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_U55 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n247), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n246), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n261) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_U54 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n245), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n260), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n244), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n243), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n249) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_U53 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n242), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n260) );
  NOR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_U52 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n241), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n240), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n239), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n251) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_U51 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n263), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n252) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_U50 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n247), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n246), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n263) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_U49 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n265), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n238), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n246) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_U48 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n244), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n238), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n254) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_U47 ( .A(
        Red_StateRegOutput[91]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n237), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n278) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_U46 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n238), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n236), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n235), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n237) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_U45 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n238), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n234), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n233), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n235) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_U44 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n244), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n247), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n259), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n248), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n233) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_U43 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n232), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n264), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n239), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n255), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n236) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_U42 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n257), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n241), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n255) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_U41 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n257), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n265), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n242), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n231), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n232) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_U40 ( .A(
        Red_StateRegOutput[93]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n230), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n279) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_U39 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n229), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n259), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n228), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n257), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n227), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n230) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_U38 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n226), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n225), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n224), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n223), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n227) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_U37 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n257), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n244), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n223) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_U36 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n222), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n224) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_U35 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n241), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n266), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n225) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_U34 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n257), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n239), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n266) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_U33 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n242), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n248), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n239) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_U32 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n259), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n257) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_U31 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n234), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n221), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n228) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_U30 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n222), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n247), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n231), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n240), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n221) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_U29 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n241), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n248), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n231) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_U28 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n273), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n248) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_U27 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n273), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n238), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n222) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_U26 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n273), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n245), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n244), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n247), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n234) );
  AND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_U25 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n270), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n264), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n247) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_U24 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n265), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n242), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n244) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_U23 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n240), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n265) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_U22 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n240), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n270), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n245) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_U21 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n241), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n270) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_U20 ( .A(
        Red_StateRegOutput[96]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n220), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n273) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_U19 ( .A(
        F_SD2_RedSB_inst_n71), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n219), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n259) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_U18 ( .A(
        Red_StateRegOutput[93]), .B(F_SD2_RedSB_inst_n69), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n219) );
  NOR4_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_U17 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n242), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n241), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n240), .A4(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n269), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n229) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_U16 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n243), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n269) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_U15 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n264), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n226), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n243) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_U14 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n238), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n226) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_U13 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n218), .B(
        Red_StateRegOutput[91]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n238) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_U12 ( .A(
        F_SD2_RedSB_inst_n69), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n217), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n218) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_U11 ( .A(
        Red_StateRegOutput[95]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n217), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n264) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_U10 ( .A(
        F_SD2_RedSB_inst_n71), .B(F_SD2_RedSB_inst_n70), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n217) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_U9 ( .A(
        Red_StateRegOutput[97]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n216), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n240) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_U8 ( .A(
        F_SD2_RedSB_inst_n71), .B(F_SD2_RedSB_inst_n72), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n216) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_U7 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n215), .B(
        Red_StateRegOutput[94]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n241) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_U6 ( .A(
        F_SD2_RedSB_inst_n69), .B(F_SD2_RedSB_inst_n72), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n215) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_U5 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n214), .B(
        Red_StateRegOutput[92]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n242) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_U4 ( .A(
        F_SD2_RedSB_inst_n69), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n220), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n214) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_U3 ( .A(
        F_SD2_RedSB_inst_n70), .B(F_SD2_RedSB_inst_n72), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_92_n220) );
  MUX2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_U54 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n240), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n239), .S(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n238), .Z(Red_Feedback[16])
         );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_U53 ( .A(
        Red_StateRegOutput[93]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n237), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n238) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_U52 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n236), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n235), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n234), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n233), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n237) );
  OR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_U51 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n232), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n231), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n230), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n233) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_U50 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n229), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n228), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n227), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n234) );
  AOI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_U49 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n226), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n225), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n224), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n223), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n236) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_U48 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n222), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n221), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n220), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n221), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n219), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n223) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_U47 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n226), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n225), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n218), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n221) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_U46 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n217), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n216), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n225) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_U45 ( .A(
        Red_StateRegOutput[96]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n215), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n239) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_U44 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n214), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n230), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n213), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n212), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n215) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_U43 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n228), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n226), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n211), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n232), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n212) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_U42 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n210), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n228), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n210), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n226), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n216), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n213) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_U41 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n220), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n216) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_U40 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n209), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n226) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_U39 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n208), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n207), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n228) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_U38 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n219), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n206), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n205), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n210) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_U37 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n219), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n206), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n208), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n205) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_U36 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n235), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n208) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_U35 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n222), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n204), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n229), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n214) );
  AND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_U34 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n206), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n219), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n204) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_U33 ( .A(
        Red_StateRegOutput[92]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n203), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n240) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_U32 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n202), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n201), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n200), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n201), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n199), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n203) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_U31 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n198), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n197), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n230), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n209), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n199) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_U30 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n227), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n220), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n218), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n197) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_U29 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n207), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n218) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_U28 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n222), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n201), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n227) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_U27 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n198), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n230), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n209), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n230), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n217), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n200) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_U26 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n231), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n206), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n209) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_U25 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n207), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n235), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n220), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n230) );
  AOI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_U24 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n229), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n211), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n207), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n224), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n198) );
  NOR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_U23 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n231), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n220), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n201), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n224) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_U22 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n219), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n220), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n211) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_U21 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n196), .B(
        Red_StateRegOutput[96]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n220) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_U20 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n201), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n219) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_U19 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n232), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n206), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n229) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_U18 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n195), .B(
        Red_StateRegOutput[95]), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n206) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_U17 ( .A(
        F_SD2_RedSB_inst_n71), .B(F_SD2_RedSB_inst_n70), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n195) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_U16 ( .A(
        Red_StateRegOutput[97]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n194), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n201) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_U15 ( .A(
        F_SD2_RedSB_inst_n71), .B(F_SD2_RedSB_inst_n72), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n194) );
  NOR4_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_U14 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n207), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n231), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n232), .A4(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n235), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n202) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_U13 ( .A(
        Red_StateRegOutput[93]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n193), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n235) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_U12 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n217), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n232) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_U11 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n192), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n193), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n217) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_U10 ( .A(
        F_SD2_RedSB_inst_n69), .B(F_SD2_RedSB_inst_n71), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n193) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_U9 ( .A(
        F_SD2_RedSB_inst_n70), .B(Red_StateRegOutput[91]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n192) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_U8 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n222), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n231) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_U7 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n191), .B(
        Red_StateRegOutput[94]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n222) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_U6 ( .A(
        F_SD2_RedSB_inst_n69), .B(F_SD2_RedSB_inst_n72), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n191) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_U5 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n190), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n196), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n207) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_U4 ( .A(
        F_SD2_RedSB_inst_n70), .B(F_SD2_RedSB_inst_n72), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n196) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_U3 ( .A(
        F_SD2_RedSB_inst_n69), .B(Red_StateRegOutput[92]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_93_n190) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_U70 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n290), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n289), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n288), .ZN(Red_Feedback[17])
         );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_U69 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n290), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n287), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n288) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_U68 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n286), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n285), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n284), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n287) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_U67 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n283), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n282), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n286), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n284) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_U66 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n289), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n285) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_U65 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n283), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n282), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n281), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n289) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_U64 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n282), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n286), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n283), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n281) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_U63 ( .A(
        Red_StateRegOutput[96]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n268), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n282) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_U62 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n267), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n266), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n265), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n269), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n268) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_U61 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n264), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n274), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n263), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n262), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n261), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n265) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_U60 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n260), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n259), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n278), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n258), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n263) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_U59 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n262), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n274) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_U58 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n273), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n272), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n264) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_U57 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n257), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n266) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_U56 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n256), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n255), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n254), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n267) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_U55 ( .A(
        Red_StateRegOutput[93]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n253), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n283) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_U54 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n252), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n262), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n251), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n250), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n253) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_U53 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n278), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n257), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n249), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n250) );
  NAND4_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_U52 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n254), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n248), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n276), .A4(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n262), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n251) );
  AOI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_U51 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n271), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n247), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n246), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n277), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n252) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_U50 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n258), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n259), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n245), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n277) );
  NOR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_U49 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n278), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n244), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n280), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n246) );
  AND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_U48 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n258), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n259), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n280) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_U47 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n243), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n259) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_U46 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n249), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n269), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n271) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_U45 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n276), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n279), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n257) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_U44 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n262), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n269), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n279) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_U43 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n244), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n256), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n245) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_U42 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n241), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n247), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n256) );
  AND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_U41 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n243), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n242), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n261) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_U40 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n278), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n272), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n242) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_U39 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n249), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n273), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n243) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_U38 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n255), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n273) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_U37 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n249), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n247), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n248) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_U36 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n275), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n255), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n254) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_U35 ( .A(
        Red_StateRegOutput[95]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n240), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n255) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_U34 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n278), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n275) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_U33 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n269), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n244) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_U32 ( .A(
        Red_StateRegOutput[96]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n239), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n269) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_U31 ( .A(
        F_SD2_RedSB_inst_n70), .B(F_SD2_RedSB_inst_n72), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n239) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_U30 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n262), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n241), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n270) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_U29 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n249), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n241) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_U28 ( .A(
        Red_StateRegOutput[94]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n238), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n249) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_U27 ( .A(
        F_SD2_RedSB_inst_n69), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n237), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n262) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_U26 ( .A(
        Red_StateRegOutput[93]), .B(F_SD2_RedSB_inst_n71), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n237) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_U25 ( .A(
        F_SD2_RedSB_inst_n70), .B(F_SD2_RedSB_inst_n71), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n240) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_U24 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n276), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n247), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n258) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_U23 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n272), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n247) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_U22 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n236), .B(
        Red_StateRegOutput[97]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n272) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_U21 ( .A(
        F_SD2_RedSB_inst_n71), .B(F_SD2_RedSB_inst_n72), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n236) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_U20 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n260), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n276) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_U19 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n235), .B(
        Red_StateRegOutput[92]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n260) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_U18 ( .A(
        F_SD2_RedSB_inst_n70), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n238), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n235) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_U17 ( .A(
        F_SD2_RedSB_inst_n69), .B(F_SD2_RedSB_inst_n72), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n238) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_U16 ( .A(
        Red_StateRegOutput[91]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n234), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n278) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_U15 ( .A(
        F_SD2_RedSB_inst_n69), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n240), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n234) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_U14 ( .A(
        Red_StateRegOutput[92]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n233), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n290) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_U13 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n258), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n229), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n231), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n232), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n233) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_U12 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n261), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n269), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n261), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n248), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n260), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n232) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_U11 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n243), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n257), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n242), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n257), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n230), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n231) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_U10 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n260), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n245), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n230) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_U9 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n278), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n270), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n244), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n254), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n229) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_U8 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n228), .B(
        Red_StateRegOutput[91]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n286) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_U7 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n224), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n277), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n227), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n228) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_U6 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n276), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n225), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n275), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n226), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n227) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_U5 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n274), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n272), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n273), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n226) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_U4 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n269), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n270), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n273), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n271), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n225) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_U3 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n280), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n279), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n278), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_94_n224) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_U73 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n281), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n280), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n281), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n279), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n278), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n282) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_U72 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n277), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n276), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n275), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n283) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_U71 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n274), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n273), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n276), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n275) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_U70 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n272), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n271), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n270), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n274) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_U69 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n269), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n276) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_U68 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n263), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n262), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n261), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n264) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_U67 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n262), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n266) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_U66 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n277), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n260) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_U65 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n258), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n257), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n277) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_U64 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n261), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n278), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n255), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n273) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_U63 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n280), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n272), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n256) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_U62 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n261), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n254), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n280) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_U61 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n271), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n279), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n262), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n251), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n252) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_U60 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n258), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n259), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n250), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n284), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n251) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_U59 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n269), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n249), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n284) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_U58 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n267), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n248), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n279) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_U57 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n285), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n271) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_U56 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n254), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n247), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n285) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_U55 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n246), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n245), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n244), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n253) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_U54 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n257), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n268), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n246), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n244) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_U53 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n270), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n243), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n242), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n245) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_U52 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n281), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n242) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_U51 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n267), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n248), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n281) );
  OR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_U50 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n272), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n249), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n248) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_U49 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n263), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n267) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_U48 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n250), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n272), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n243) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_U47 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n278), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n250) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_U46 ( .A(
        Red_StateRegOutput[91]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n241), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n286) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_U45 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n269), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n240), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n239), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n241) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_U44 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n257), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n259), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n238), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n237), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n239) );
  OR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_U43 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n246), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n268), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n265), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n237) );
  OR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_U42 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n278), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n249), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n258), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n265) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_U41 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n254), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n246) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_U40 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n263), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n247), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n262), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n236), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n249), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n238) );
  AND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_U39 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n263), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n247), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n236) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_U38 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n272), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n254), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n262) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_U37 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n261), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n278), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n247) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_U36 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n258), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n261) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_U35 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n269), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n270), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n263) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_U34 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n270), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n249), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n259) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_U33 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n268), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n270) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_U32 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n272), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n278), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n257) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_U31 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n255), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n272) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_U30 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n255), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n235), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n258), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n235), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n249), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n240) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_U29 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n234), .B(
        Red_StateRegOutput[91]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n249) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_U28 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n233), .B(
        F_SD2_RedSB_inst_n70), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n234) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_U27 ( .A(
        Red_StateRegOutput[93]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n233), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n258) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_U26 ( .A(
        F_SD2_RedSB_inst_n71), .B(F_SD2_RedSB_inst_n69), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n233) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_U25 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n254), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n278), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n268), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n235) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_U24 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n232), .B(
        Red_StateRegOutput[94]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n268) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_U23 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n231), .B(
        F_SD2_RedSB_inst_n70), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n278) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_U22 ( .A(
        Red_StateRegOutput[96]), .B(F_SD2_RedSB_inst_n72), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n231) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_U21 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n230), .B(
        Red_StateRegOutput[92]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n254) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_U20 ( .A(
        F_SD2_RedSB_inst_n70), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n232), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n230) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_U19 ( .A(
        F_SD2_RedSB_inst_n69), .B(F_SD2_RedSB_inst_n72), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n232) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_U18 ( .A(
        Red_StateRegOutput[97]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n229), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n255) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_U17 ( .A(
        F_SD2_RedSB_inst_n71), .B(F_SD2_RedSB_inst_n72), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n229) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_U16 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n228), .B(
        Red_StateRegOutput[95]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n269) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_U15 ( .A(
        F_SD2_RedSB_inst_n71), .B(F_SD2_RedSB_inst_n70), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n228) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_U14 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n286), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n218), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n226), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n224), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n227), .ZN(Red_Feedback[18])
         );
  NOR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_U13 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n218), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n224), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n226), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n227) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_U12 ( .A(
        Red_StateRegOutput[96]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n225), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n226) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_U11 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n285), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n284), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n283), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n282), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n225) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_U10 ( .B1(
        Red_StateRegOutput[93]), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n222), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n223), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n224) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_U9 ( .B1(
        Red_StateRegOutput[93]), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n222), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n286), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n223) );
  AOI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_U8 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n268), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n219), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n220), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n221), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n222) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_U7 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n285), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n259), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n260), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n268), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n221) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_U6 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n264), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n265), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n266), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n267), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n220) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_U5 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n284), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n256), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n273), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n219) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_U4 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n217), .B(
        Red_StateRegOutput[92]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n218) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_U3 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n253), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n252), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_95_n217) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_U72 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n283), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n282), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n281), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n280), .ZN(Red_Feedback[19])
         );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_U71 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n279), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n280), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n278), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n282) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_U70 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n279), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n280), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n281), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n278) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_U69 ( .A(
        Red_StateRegOutput[96]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n277), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n281) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_U68 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n276), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n275), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n277) );
  NAND4_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_U67 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n274), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n273), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n272), .A4(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n271), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n275) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_U66 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n270), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n269), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n268), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n267), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n276) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_U65 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n266), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n267) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_U64 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n273), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n265), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n264), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n263), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n269) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_U63 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n262), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n264) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_U62 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n261), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n271), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n260), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n259), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n265) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_U61 ( .A(
        Red_StateRegOutput[92]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n258), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n280) );
  NOR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_U60 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n257), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n256), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n255), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n258) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_U59 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n253), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n252), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n262) );
  AOI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_U58 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n274), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n251), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n250), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n249), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n256) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_U57 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n248), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n247), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n274), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n249) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_U56 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n270), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n246), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n251) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_U55 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n247), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n270) );
  NOR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_U54 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n253), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n246), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n252), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n257) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_U53 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n259), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n250), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n252) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_U52 ( .A(
        Red_StateRegOutput[91]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n245), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n279) );
  AOI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_U51 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n274), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n244), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n243), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n242), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n245) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_U50 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n253), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n241), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n254), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n240), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n242) );
  OR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_U49 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n253), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n241), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n259), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n240) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_U48 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n239), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n250), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n246), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n254) );
  NOR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_U47 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n239), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n238), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n271), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n243) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_U46 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n273), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n261), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n248), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n237), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n238) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_U45 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n236), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n259), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n235), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n244) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_U44 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n234), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n248), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n261), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n235) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_U43 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n233), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n236) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_U42 ( .A(
        Red_StateRegOutput[93]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n232), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n283) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_U41 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n261), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n231), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n230), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n232) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_U40 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n266), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n229), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n228), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n263), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n230) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_U39 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n246), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n227), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n263) );
  NAND4_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_U38 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n239), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n268), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n273), .A4(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n229), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n228) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_U37 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n271), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n268) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_U36 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n239), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n272), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n261), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n233), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n266) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_U35 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n247), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n250), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n233) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_U34 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n246), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n241), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n272) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_U33 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n247), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n227), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n241) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_U32 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n259), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n239) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_U31 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n273), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n226), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n225), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n253), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n231) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_U30 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n234), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n246), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n260), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n246), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n237), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n226) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_U29 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n274), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n247), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n237) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_U28 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n229), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n274) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_U27 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n253), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n260) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_U26 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n229), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n271), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n253) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_U25 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n224), .B(
        Red_StateRegOutput[95]), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n271) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_U24 ( .A(
        F_SD2_RedSB_inst_n70), .B(F_SD2_RedSB_inst_n71), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n224) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_U23 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n223), .B(
        Red_StateRegOutput[94]), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n229) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_U22 ( .A(
        F_SD2_RedSB_inst_n69), .B(F_SD2_RedSB_inst_n72), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n223) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_U21 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n248), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n246) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_U20 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n222), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n221), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n248) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_U19 ( .A(
        F_SD2_RedSB_inst_n72), .B(Red_StateRegOutput[92]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n222) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_U18 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n225), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n234) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_U17 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n259), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n247), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n225) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_U16 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n220), .B(
        Red_StateRegOutput[96]), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n247) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_U15 ( .A(
        F_SD2_RedSB_inst_n70), .B(F_SD2_RedSB_inst_n72), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n220) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_U14 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n219), .B(
        F_SD2_RedSB_inst_n71), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n259) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_U13 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n221), .B(
        Red_StateRegOutput[91]), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n219) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_U12 ( .A(
        F_SD2_RedSB_inst_n69), .B(F_SD2_RedSB_inst_n70), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n221) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_U11 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n250), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n273) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_U10 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n218), .B(
        Red_StateRegOutput[97]), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n250) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_U9 ( .A(
        F_SD2_RedSB_inst_n71), .B(F_SD2_RedSB_inst_n72), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n218) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_U8 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n227), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n261) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_U7 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n217), .B(
        F_SD2_RedSB_inst_n71), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n227) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_U6 ( .A(
        Red_StateRegOutput[93]), .B(F_SD2_RedSB_inst_n69), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n217) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_U5 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n254), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n215), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n216), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n255) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_U4 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n272), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n262), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n216) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_U3 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n268), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n270), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n261), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n274), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_96_n215) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_U65 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n283), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n282), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n281), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n280), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n279), .ZN(Red_Feedback[20])
         );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_U64 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n283), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n282), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n281), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n279) );
  MUX2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_U63 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n283), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n282), .S(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n278), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n280) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_U62 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n277), .B(
        Red_StateRegOutput[93]), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n278) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_U61 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n276), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n275), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n274), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n277) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_U60 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n273), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n274) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_U59 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n272), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n271), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n270), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n269), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n268), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n273) );
  AND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_U58 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n267), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n266), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n265), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n269) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_U57 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n266), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n264), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n263), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n262), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n275) );
  AOI222_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_U56 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n261), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n260), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n261), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n259), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n260), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n259), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n263) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_U55 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n258), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n268), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n259) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_U54 ( .A(
        Red_StateRegOutput[91]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n257), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n281) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_U53 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n268), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n256), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n255), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n257) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_U52 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n268), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n254), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n262), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n255) );
  AOI222_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_U51 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n261), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n260), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n261), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n253), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n260), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n253), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n254) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_U50 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n276), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n258), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n253) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_U49 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n252), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n251), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n250), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n249), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n256) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_U48 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n276), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n266), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n248), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n247), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n252) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_U47 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n264), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n247) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_U46 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n272), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n258), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n264) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_U45 ( .A(
        Red_StateRegOutput[92]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n246), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n282) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_U44 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n248), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n262), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n245), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n244), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n246) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_U43 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n248), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n243), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n244) );
  AOI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_U42 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n271), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n242), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n241), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n240), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n245) );
  NOR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_U41 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n270), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n239), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n250), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n240) );
  AND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_U40 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n238), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n268), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n260), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n241) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_U39 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n248), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n266), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n260) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_U38 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n251), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n237), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n249), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n238) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_U37 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n276), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n270), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n249) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_U36 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n258), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n236), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n262) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_U35 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n237), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n258) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_U34 ( .A(
        Red_StateRegOutput[96]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n235), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n283) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_U33 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n234), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n237), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n233), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n237), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n232), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n235) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_U32 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n251), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n268), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n267), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n236), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n271), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n232) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_U31 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n250), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n276), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n271) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_U30 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n237), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n248), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n250) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_U29 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n239), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n272), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n236) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_U28 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n242), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n265), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n243), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n233) );
  AND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_U27 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n261), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n231), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n243) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_U26 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n276), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n248), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n265) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_U25 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n230), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n229), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n248) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_U24 ( .A(
        F_SD2_RedSB_inst_n69), .B(Red_StateRegOutput[92]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n230) );
  OR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_U23 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n261), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n231), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n242) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_U22 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n268), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n266), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n231) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_U21 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n228), .B(
        Red_StateRegOutput[91]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n268) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_U20 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n227), .B(
        F_SD2_RedSB_inst_n70), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n228) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_U19 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n267), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n270), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n261) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_U18 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n272), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n270) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_U17 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n226), .B(
        Red_StateRegOutput[94]), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n272) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_U16 ( .A(
        F_SD2_RedSB_inst_n69), .B(F_SD2_RedSB_inst_n72), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n226) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_U15 ( .A(
        Red_StateRegOutput[96]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n229), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n237) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_U14 ( .A(
        F_SD2_RedSB_inst_n72), .B(F_SD2_RedSB_inst_n70), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n229) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_U13 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n225), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n234) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_U12 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n267), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n239), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n224), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n225) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_U11 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n267), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n239), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n276), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n224) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_U10 ( .A(
        Red_StateRegOutput[93]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n227), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n276) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_U9 ( .A(
        F_SD2_RedSB_inst_n71), .B(F_SD2_RedSB_inst_n69), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n227) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_U8 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n266), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n239) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_U7 ( .A(
        Red_StateRegOutput[97]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n223), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n266) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_U6 ( .A(
        F_SD2_RedSB_inst_n71), .B(F_SD2_RedSB_inst_n72), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n223) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_U5 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n251), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n267) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_U4 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n222), .B(
        Red_StateRegOutput[95]), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n251) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_U3 ( .A(
        F_SD2_RedSB_inst_n71), .B(F_SD2_RedSB_inst_n70), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_97_n222) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_U69 ( .A(
        Red_StateRegOutput[99]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n280), .Z(Red_Feedback[21])
         );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_U68 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n279), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n278), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n280) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_U67 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n277), .B2(
        Red_StateRegOutput[100]), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n276), .C2(
        Red_StateRegOutput[103]), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n275), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n278) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_U66 ( .A1(
        Red_StateRegOutput[100]), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n277), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n276), .B2(
        Red_StateRegOutput[103]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n275) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_U65 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n274), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n273), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n276) );
  AOI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_U64 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n272), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n271), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n270), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n269), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n273) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_U63 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n268), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n267), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n266), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n265), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n264), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n269) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_U62 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n268), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n263), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n262), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n270) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_U61 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n268), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n263), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n261), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n262) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_U60 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n260), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n259), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n258), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n271) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_U59 ( .A(
        Red_StateRegOutput[98]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n257), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n274) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_U58 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n253), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n252), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n251), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n254) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_U57 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n252), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n253), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n250), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n255) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_U56 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n245), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n244), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n243), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n242), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n249) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_U55 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n241), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n240), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n242), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n239), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n238), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n277) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_U54 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n237), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n236), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n235), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n238) );
  AOI222_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_U53 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n253), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n251), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n253), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n234), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n251), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n234), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n236) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_U52 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n244), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n267), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n234) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_U51 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n263), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n248), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n251) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_U50 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n233), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n253) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_U49 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n256), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n232), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n239) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_U48 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n261), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n263), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n231), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n240) );
  NOR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_U47 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n267), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n246), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n259), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n231) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_U46 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n247), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n248), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n259) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_U45 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n268), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n230), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n246) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_U44 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n256), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n267) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_U43 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n244), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n247), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n261) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_U42 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n264), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n260), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n229), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n279) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_U41 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n248), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n228), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n227), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n229) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_U40 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n248), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n226), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n250), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n227) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_U39 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n237), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n250) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_U38 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n244), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n265), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n237) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_U37 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n241), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n230), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n265) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_U36 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n243), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n245), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n256), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n263), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n226) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_U35 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n242), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n247), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n245) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_U34 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n266), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n244), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n243) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_U33 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n272), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n225), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n258), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n228) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_U32 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n233), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n224), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n258) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_U31 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n242), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n230), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n225) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_U30 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n233), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n224), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n260) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_U29 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n230), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n256), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n224) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_U28 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n223), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n222), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n256) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_U27 ( .A(
        Red_StateRegOutput[98]), .B(F_SD2_RedSB_inst_n73), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n223) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_U26 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n263), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n230) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_U25 ( .A(
        Red_StateRegOutput[104]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n221), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n263) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_U24 ( .A(
        F_SD2_RedSB_inst_n76), .B(F_SD2_RedSB_inst_n75), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n221) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_U23 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n241), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n268), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n233) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_U22 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n266), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n268) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_U21 ( .A(
        Red_StateRegOutput[102]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n222), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n266) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_U20 ( .A(
        F_SD2_RedSB_inst_n74), .B(F_SD2_RedSB_inst_n75), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n222) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_U19 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n242), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n241) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_U18 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n220), .B(
        Red_StateRegOutput[101]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n242) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_U17 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n232), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n264) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_U16 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n252), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n248), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n232) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_U15 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n219), .B(
        F_SD2_RedSB_inst_n74), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n248) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_U14 ( .A(
        Red_StateRegOutput[99]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n220), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n219) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_U13 ( .A(
        F_SD2_RedSB_inst_n76), .B(F_SD2_RedSB_inst_n73), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n220) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_U12 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n244), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n247), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n252) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_U11 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n235), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n247) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_U10 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n218), .B(
        Red_StateRegOutput[100]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n235) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_U9 ( .A(
        F_SD2_RedSB_inst_n73), .B(F_SD2_RedSB_inst_n75), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n218) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_U8 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n272), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n244) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_U7 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n217), .B(
        F_SD2_RedSB_inst_n74), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n272) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_U6 ( .A(
        Red_StateRegOutput[103]), .B(F_SD2_RedSB_inst_n76), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n217) );
  OAI33_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_U5 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n256), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n215), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n216), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n267), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n255), .B3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n254), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n257) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_U4 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n249), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n248), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n216) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_U3 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n247), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n246), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_98_n215) );
  AOI222_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_U69 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n279), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n278), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n279), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n277), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n278), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n276), .ZN(Red_Feedback[22])
         );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_U68 ( .A(
        Red_StateRegOutput[103]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n275), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n276) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_U67 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n274), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n273), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n272), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n273), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n271), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n275) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_U66 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n270), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n269), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n268), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n269), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n267), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n271) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_U65 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n266), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n267) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_U64 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n265), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n264), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n268) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_U63 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n263), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n262), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n261), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n272) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_U62 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n260), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n259), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n262) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_U61 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n265), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n264), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n258), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n274) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_U60 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n265), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n264), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n257), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n258) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_U59 ( .A(
        Red_StateRegOutput[99]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n256), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n277) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_U58 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n255), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n254), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n253), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n256) );
  AOI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_U57 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n266), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n252), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n251), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n250), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n253) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_U56 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n249), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n248), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n260), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n261), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n250) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_U55 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n247), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n246), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n261) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_U54 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n245), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n260), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n244), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n243), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n249) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_U53 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n242), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n260) );
  NOR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_U52 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n241), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n240), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n239), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n251) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_U51 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n263), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n252) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_U50 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n247), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n246), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n263) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_U49 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n265), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n238), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n246) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_U48 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n244), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n238), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n254) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_U47 ( .A(
        Red_StateRegOutput[98]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n237), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n278) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_U46 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n238), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n236), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n235), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n237) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_U45 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n238), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n234), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n233), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n235) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_U44 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n244), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n247), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n259), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n248), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n233) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_U43 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n232), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n264), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n239), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n255), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n236) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_U42 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n257), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n241), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n255) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_U41 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n257), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n265), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n242), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n231), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n232) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_U40 ( .A(
        Red_StateRegOutput[100]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n230), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n279) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_U39 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n229), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n259), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n228), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n257), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n227), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n230) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_U38 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n226), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n225), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n224), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n223), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n227) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_U37 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n257), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n244), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n223) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_U36 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n222), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n224) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_U35 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n241), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n266), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n225) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_U34 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n257), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n239), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n266) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_U33 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n242), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n248), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n239) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_U32 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n259), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n257) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_U31 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n234), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n221), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n228) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_U30 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n222), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n247), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n231), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n240), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n221) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_U29 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n241), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n248), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n231) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_U28 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n273), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n248) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_U27 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n273), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n238), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n222) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_U26 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n273), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n245), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n244), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n247), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n234) );
  AND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_U25 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n270), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n264), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n247) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_U24 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n265), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n242), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n244) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_U23 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n240), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n265) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_U22 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n240), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n270), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n245) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_U21 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n241), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n270) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_U20 ( .A(
        Red_StateRegOutput[103]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n220), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n273) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_U19 ( .A(
        F_SD2_RedSB_inst_n75), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n219), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n259) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_U18 ( .A(
        Red_StateRegOutput[100]), .B(F_SD2_RedSB_inst_n73), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n219) );
  NOR4_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_U17 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n242), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n241), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n240), .A4(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n269), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n229) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_U16 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n243), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n269) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_U15 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n264), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n226), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n243) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_U14 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n238), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n226) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_U13 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n218), .B(
        Red_StateRegOutput[98]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n238) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_U12 ( .A(
        F_SD2_RedSB_inst_n73), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n217), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n218) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_U11 ( .A(
        Red_StateRegOutput[102]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n217), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n264) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_U10 ( .A(
        F_SD2_RedSB_inst_n75), .B(F_SD2_RedSB_inst_n74), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n217) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_U9 ( .A(
        Red_StateRegOutput[104]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n216), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n240) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_U8 ( .A(
        F_SD2_RedSB_inst_n75), .B(F_SD2_RedSB_inst_n76), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n216) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_U7 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n215), .B(
        Red_StateRegOutput[101]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n241) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_U6 ( .A(
        F_SD2_RedSB_inst_n73), .B(F_SD2_RedSB_inst_n76), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n215) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_U5 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n214), .B(
        Red_StateRegOutput[99]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n242) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_U4 ( .A(
        F_SD2_RedSB_inst_n73), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n220), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n214) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_U3 ( .A(
        F_SD2_RedSB_inst_n74), .B(F_SD2_RedSB_inst_n76), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_99_n220) );
  MUX2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_U54 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n240), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n239), .S(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n238), .Z(Red_Feedback[23])
         );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_U53 ( .A(
        Red_StateRegOutput[100]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n237), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n238) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_U52 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n236), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n235), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n234), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n233), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n237) );
  OR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_U51 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n232), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n231), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n230), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n233) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_U50 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n229), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n228), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n227), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n234) );
  AOI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_U49 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n226), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n225), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n224), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n223), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n236) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_U48 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n222), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n221), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n220), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n221), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n219), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n223) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_U47 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n226), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n225), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n218), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n221) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_U46 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n217), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n216), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n225) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_U45 ( .A(
        Red_StateRegOutput[103]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n215), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n239) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_U44 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n214), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n230), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n213), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n212), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n215) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_U43 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n228), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n226), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n211), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n232), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n212) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_U42 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n210), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n228), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n210), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n226), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n216), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n213) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_U41 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n220), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n216) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_U40 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n209), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n226) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_U39 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n208), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n207), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n228) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_U38 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n219), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n206), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n205), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n210) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_U37 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n219), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n206), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n208), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n205) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_U36 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n235), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n208) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_U35 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n222), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n204), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n229), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n214) );
  AND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_U34 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n206), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n219), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n204) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_U33 ( .A(
        Red_StateRegOutput[99]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n203), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n240) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_U32 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n202), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n201), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n200), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n201), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n199), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n203) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_U31 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n198), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n197), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n230), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n209), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n199) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_U30 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n227), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n220), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n218), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n197) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_U29 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n207), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n218) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_U28 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n222), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n201), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n227) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_U27 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n198), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n230), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n209), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n230), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n217), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n200) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_U26 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n231), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n206), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n209) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_U25 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n207), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n235), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n220), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n230) );
  AOI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_U24 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n229), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n211), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n207), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n224), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n198) );
  NOR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_U23 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n231), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n220), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n201), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n224) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_U22 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n219), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n220), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n211) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_U21 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n196), .B(
        Red_StateRegOutput[103]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n220) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_U20 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n201), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n219) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_U19 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n232), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n206), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n229) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_U18 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n195), .B(
        Red_StateRegOutput[102]), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n206) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_U17 ( .A(
        F_SD2_RedSB_inst_n75), .B(F_SD2_RedSB_inst_n74), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n195) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_U16 ( .A(
        Red_StateRegOutput[104]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n194), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n201) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_U15 ( .A(
        F_SD2_RedSB_inst_n75), .B(F_SD2_RedSB_inst_n76), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n194) );
  NOR4_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_U14 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n207), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n231), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n232), .A4(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n235), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n202) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_U13 ( .A(
        Red_StateRegOutput[100]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n193), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n235) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_U12 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n217), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n232) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_U11 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n192), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n193), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n217) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_U10 ( .A(
        F_SD2_RedSB_inst_n73), .B(F_SD2_RedSB_inst_n75), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n193) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_U9 ( .A(
        F_SD2_RedSB_inst_n74), .B(Red_StateRegOutput[98]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n192) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_U8 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n222), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n231) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_U7 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n191), .B(
        Red_StateRegOutput[101]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n222) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_U6 ( .A(
        F_SD2_RedSB_inst_n73), .B(F_SD2_RedSB_inst_n76), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n191) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_U5 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n190), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n196), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n207) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_U4 ( .A(
        F_SD2_RedSB_inst_n74), .B(F_SD2_RedSB_inst_n76), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n196) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_U3 ( .A(
        F_SD2_RedSB_inst_n73), .B(Red_StateRegOutput[99]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_100_n190) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_U70 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n290), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n289), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n288), .ZN(Red_Feedback[24])
         );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_U69 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n290), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n287), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n288) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_U68 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n286), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n285), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n284), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n287) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_U67 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n283), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n282), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n286), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n284) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_U66 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n289), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n285) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_U65 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n283), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n282), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n281), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n289) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_U64 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n282), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n286), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n283), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n281) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_U63 ( .A(
        Red_StateRegOutput[103]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n268), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n282) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_U62 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n267), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n266), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n265), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n269), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n268) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_U61 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n264), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n274), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n263), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n262), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n261), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n265) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_U60 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n260), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n259), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n278), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n258), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n263) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_U59 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n262), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n274) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_U58 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n273), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n272), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n264) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_U57 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n257), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n266) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_U56 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n256), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n255), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n254), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n267) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_U55 ( .A(
        Red_StateRegOutput[100]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n253), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n283) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_U54 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n252), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n262), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n251), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n250), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n253) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_U53 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n278), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n257), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n249), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n250) );
  NAND4_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_U52 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n254), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n248), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n276), .A4(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n262), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n251) );
  AOI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_U51 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n271), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n247), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n246), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n277), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n252) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_U50 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n258), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n259), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n245), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n277) );
  NOR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_U49 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n278), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n244), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n280), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n246) );
  AND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_U48 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n258), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n259), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n280) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_U47 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n243), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n259) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_U46 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n249), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n269), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n271) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_U45 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n276), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n279), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n257) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_U44 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n262), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n269), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n279) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_U43 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n244), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n256), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n245) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_U42 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n241), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n247), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n256) );
  AND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_U41 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n243), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n242), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n261) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_U40 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n278), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n272), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n242) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_U39 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n249), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n273), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n243) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_U38 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n255), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n273) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_U37 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n249), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n247), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n248) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_U36 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n275), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n255), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n254) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_U35 ( .A(
        Red_StateRegOutput[102]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n240), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n255) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_U34 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n278), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n275) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_U33 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n269), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n244) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_U32 ( .A(
        Red_StateRegOutput[103]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n239), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n269) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_U31 ( .A(
        F_SD2_RedSB_inst_n74), .B(F_SD2_RedSB_inst_n76), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n239) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_U30 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n262), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n241), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n270) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_U29 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n249), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n241) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_U28 ( .A(
        Red_StateRegOutput[101]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n238), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n249) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_U27 ( .A(
        F_SD2_RedSB_inst_n73), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n237), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n262) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_U26 ( .A(
        Red_StateRegOutput[100]), .B(F_SD2_RedSB_inst_n75), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n237) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_U25 ( .A(
        F_SD2_RedSB_inst_n74), .B(F_SD2_RedSB_inst_n75), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n240) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_U24 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n276), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n247), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n258) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_U23 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n272), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n247) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_U22 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n236), .B(
        Red_StateRegOutput[104]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n272) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_U21 ( .A(
        F_SD2_RedSB_inst_n75), .B(F_SD2_RedSB_inst_n76), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n236) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_U20 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n260), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n276) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_U19 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n235), .B(
        Red_StateRegOutput[99]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n260) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_U18 ( .A(
        F_SD2_RedSB_inst_n74), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n238), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n235) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_U17 ( .A(
        F_SD2_RedSB_inst_n73), .B(F_SD2_RedSB_inst_n76), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n238) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_U16 ( .A(
        Red_StateRegOutput[98]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n234), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n278) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_U15 ( .A(
        F_SD2_RedSB_inst_n73), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n240), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n234) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_U14 ( .A(
        Red_StateRegOutput[99]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n233), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n290) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_U13 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n258), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n229), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n231), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n232), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n233) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_U12 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n261), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n269), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n261), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n248), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n260), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n232) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_U11 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n243), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n257), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n242), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n257), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n230), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n231) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_U10 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n260), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n245), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n230) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_U9 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n278), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n270), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n244), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n254), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n229) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_U8 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n228), .B(
        Red_StateRegOutput[98]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n286) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_U7 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n224), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n277), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n227), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n228) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_U6 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n276), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n225), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n275), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n226), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n227) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_U5 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n274), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n272), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n273), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n226) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_U4 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n269), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n270), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n273), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n271), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n225) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_U3 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n280), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n279), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n278), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_101_n224) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_U73 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n281), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n280), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n281), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n279), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n278), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n282) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_U72 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n277), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n276), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n275), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n283) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_U71 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n274), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n273), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n276), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n275) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_U70 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n272), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n271), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n270), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n274) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_U69 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n269), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n276) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_U68 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n263), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n262), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n261), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n264) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_U67 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n262), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n266) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_U66 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n277), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n260) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_U65 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n258), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n257), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n277) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_U64 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n261), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n278), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n255), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n273) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_U63 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n280), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n272), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n256) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_U62 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n261), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n254), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n280) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_U61 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n271), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n279), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n262), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n251), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n252) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_U60 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n258), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n259), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n250), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n284), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n251) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_U59 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n269), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n249), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n284) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_U58 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n267), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n248), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n279) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_U57 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n285), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n271) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_U56 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n254), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n247), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n285) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_U55 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n246), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n245), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n244), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n253) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_U54 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n257), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n268), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n246), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n244) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_U53 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n270), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n243), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n242), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n245) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_U52 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n281), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n242) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_U51 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n267), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n248), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n281) );
  OR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_U50 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n272), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n249), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n248) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_U49 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n263), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n267) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_U48 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n250), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n272), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n243) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_U47 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n278), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n250) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_U46 ( .A(
        Red_StateRegOutput[98]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n241), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n286) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_U45 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n269), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n240), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n239), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n241) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_U44 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n257), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n259), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n238), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n237), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n239) );
  OR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_U43 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n246), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n268), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n265), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n237) );
  OR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_U42 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n278), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n249), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n258), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n265) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_U41 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n254), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n246) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_U40 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n263), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n247), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n262), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n236), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n249), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n238) );
  AND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_U39 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n263), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n247), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n236) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_U38 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n272), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n254), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n262) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_U37 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n261), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n278), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n247) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_U36 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n258), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n261) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_U35 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n269), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n270), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n263) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_U34 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n270), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n249), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n259) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_U33 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n268), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n270) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_U32 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n272), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n278), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n257) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_U31 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n255), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n272) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_U30 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n255), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n235), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n258), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n235), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n249), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n240) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_U29 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n234), .B(
        Red_StateRegOutput[98]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n249) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_U28 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n233), .B(
        F_SD2_RedSB_inst_n74), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n234) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_U27 ( .A(
        Red_StateRegOutput[100]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n233), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n258) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_U26 ( .A(
        F_SD2_RedSB_inst_n75), .B(F_SD2_RedSB_inst_n73), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n233) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_U25 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n254), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n278), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n268), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n235) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_U24 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n232), .B(
        Red_StateRegOutput[101]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n268) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_U23 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n231), .B(
        F_SD2_RedSB_inst_n74), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n278) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_U22 ( .A(
        Red_StateRegOutput[103]), .B(F_SD2_RedSB_inst_n76), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n231) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_U21 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n230), .B(
        Red_StateRegOutput[99]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n254) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_U20 ( .A(
        F_SD2_RedSB_inst_n74), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n232), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n230) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_U19 ( .A(
        F_SD2_RedSB_inst_n73), .B(F_SD2_RedSB_inst_n76), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n232) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_U18 ( .A(
        Red_StateRegOutput[104]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n229), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n255) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_U17 ( .A(
        F_SD2_RedSB_inst_n75), .B(F_SD2_RedSB_inst_n76), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n229) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_U16 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n228), .B(
        Red_StateRegOutput[102]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n269) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_U15 ( .A(
        F_SD2_RedSB_inst_n75), .B(F_SD2_RedSB_inst_n74), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n228) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_U14 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n286), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n218), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n226), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n224), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n227), .ZN(Red_Feedback[25])
         );
  NOR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_U13 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n218), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n224), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n226), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n227) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_U12 ( .A(
        Red_StateRegOutput[103]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n225), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n226) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_U11 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n285), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n284), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n283), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n282), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n225) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_U10 ( .B1(
        Red_StateRegOutput[100]), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n222), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n223), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n224) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_U9 ( .B1(
        Red_StateRegOutput[100]), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n222), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n286), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n223) );
  AOI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_U8 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n268), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n219), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n220), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n221), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n222) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_U7 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n285), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n259), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n260), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n268), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n221) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_U6 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n264), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n265), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n266), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n267), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n220) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_U5 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n284), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n256), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n273), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n219) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_U4 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n217), .B(
        Red_StateRegOutput[99]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n218) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_U3 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n253), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n252), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_102_n217) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_U72 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n283), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n282), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n281), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n280), .ZN(Red_Feedback[26])
         );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_U71 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n279), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n280), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n278), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n282) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_U70 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n279), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n280), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n281), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n278) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_U69 ( .A(
        Red_StateRegOutput[103]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n277), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n281) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_U68 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n276), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n275), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n277) );
  NAND4_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_U67 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n274), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n273), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n272), .A4(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n271), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n275) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_U66 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n270), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n269), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n268), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n267), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n276) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_U65 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n266), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n267) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_U64 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n273), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n265), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n264), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n263), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n269) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_U63 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n262), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n264) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_U62 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n261), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n271), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n260), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n259), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n265) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_U61 ( .A(
        Red_StateRegOutput[99]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n258), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n280) );
  NOR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_U60 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n257), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n256), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n255), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n258) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_U59 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n253), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n252), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n262) );
  AOI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_U58 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n274), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n251), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n250), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n249), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n256) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_U57 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n248), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n247), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n274), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n249) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_U56 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n270), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n246), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n251) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_U55 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n247), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n270) );
  NOR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_U54 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n253), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n246), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n252), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n257) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_U53 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n259), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n250), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n252) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_U52 ( .A(
        Red_StateRegOutput[98]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n245), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n279) );
  AOI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_U51 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n274), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n244), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n243), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n242), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n245) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_U50 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n253), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n241), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n254), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n240), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n242) );
  OR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_U49 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n253), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n241), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n259), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n240) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_U48 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n239), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n250), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n246), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n254) );
  NOR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_U47 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n239), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n238), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n271), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n243) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_U46 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n273), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n261), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n248), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n237), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n238) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_U45 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n236), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n259), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n235), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n244) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_U44 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n234), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n248), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n261), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n235) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_U43 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n233), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n236) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_U42 ( .A(
        Red_StateRegOutput[100]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n232), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n283) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_U41 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n261), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n231), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n230), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n232) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_U40 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n266), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n229), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n228), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n263), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n230) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_U39 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n246), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n227), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n263) );
  NAND4_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_U38 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n239), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n268), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n273), .A4(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n229), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n228) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_U37 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n271), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n268) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_U36 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n239), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n272), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n261), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n233), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n266) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_U35 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n247), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n250), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n233) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_U34 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n246), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n241), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n272) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_U33 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n247), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n227), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n241) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_U32 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n259), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n239) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_U31 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n273), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n226), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n225), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n253), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n231) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_U30 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n234), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n246), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n260), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n246), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n237), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n226) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_U29 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n274), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n247), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n237) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_U28 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n229), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n274) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_U27 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n253), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n260) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_U26 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n229), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n271), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n253) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_U25 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n224), .B(
        Red_StateRegOutput[102]), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n271) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_U24 ( .A(
        F_SD2_RedSB_inst_n74), .B(F_SD2_RedSB_inst_n75), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n224) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_U23 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n223), .B(
        Red_StateRegOutput[101]), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n229) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_U22 ( .A(
        F_SD2_RedSB_inst_n73), .B(F_SD2_RedSB_inst_n76), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n223) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_U21 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n248), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n246) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_U20 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n222), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n221), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n248) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_U19 ( .A(
        F_SD2_RedSB_inst_n76), .B(Red_StateRegOutput[99]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n222) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_U18 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n225), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n234) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_U17 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n259), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n247), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n225) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_U16 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n220), .B(
        Red_StateRegOutput[103]), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n247) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_U15 ( .A(
        F_SD2_RedSB_inst_n74), .B(F_SD2_RedSB_inst_n76), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n220) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_U14 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n219), .B(
        F_SD2_RedSB_inst_n75), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n259) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_U13 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n221), .B(
        Red_StateRegOutput[98]), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n219) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_U12 ( .A(
        F_SD2_RedSB_inst_n73), .B(F_SD2_RedSB_inst_n74), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n221) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_U11 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n250), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n273) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_U10 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n218), .B(
        Red_StateRegOutput[104]), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n250) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_U9 ( .A(
        F_SD2_RedSB_inst_n75), .B(F_SD2_RedSB_inst_n76), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n218) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_U8 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n227), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n261) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_U7 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n217), .B(
        F_SD2_RedSB_inst_n75), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n227) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_U6 ( .A(
        Red_StateRegOutput[100]), .B(F_SD2_RedSB_inst_n73), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n217) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_U5 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n254), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n215), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n216), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n255) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_U4 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n272), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n262), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n216) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_U3 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n268), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n270), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n261), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n274), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_103_n215) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_U65 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n283), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n282), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n281), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n280), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n279), .ZN(Red_Feedback[27])
         );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_U64 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n283), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n282), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n281), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n279) );
  MUX2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_U63 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n283), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n282), .S(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n278), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n280) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_U62 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n277), .B(
        Red_StateRegOutput[100]), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n278) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_U61 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n276), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n275), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n274), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n277) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_U60 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n273), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n274) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_U59 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n272), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n271), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n270), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n269), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n268), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n273) );
  AND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_U58 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n267), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n266), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n265), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n269) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_U57 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n266), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n264), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n263), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n262), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n275) );
  AOI222_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_U56 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n261), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n260), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n261), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n259), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n260), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n259), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n263) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_U55 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n258), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n268), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n259) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_U54 ( .A(
        Red_StateRegOutput[98]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n257), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n281) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_U53 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n268), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n256), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n255), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n257) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_U52 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n268), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n254), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n262), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n255) );
  AOI222_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_U51 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n261), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n260), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n261), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n253), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n260), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n253), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n254) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_U50 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n276), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n258), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n253) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_U49 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n252), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n251), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n250), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n249), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n256) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_U48 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n276), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n266), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n248), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n247), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n252) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_U47 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n264), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n247) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_U46 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n272), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n258), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n264) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_U45 ( .A(
        Red_StateRegOutput[99]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n246), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n282) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_U44 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n248), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n262), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n245), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n244), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n246) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_U43 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n248), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n243), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n244) );
  AOI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_U42 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n271), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n242), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n241), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n240), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n245) );
  NOR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_U41 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n270), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n239), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n250), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n240) );
  AND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_U40 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n238), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n268), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n260), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n241) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_U39 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n248), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n266), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n260) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_U38 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n251), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n237), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n249), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n238) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_U37 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n276), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n270), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n249) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_U36 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n258), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n236), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n262) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_U35 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n237), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n258) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_U34 ( .A(
        Red_StateRegOutput[103]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n235), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n283) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_U33 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n234), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n237), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n233), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n237), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n232), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n235) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_U32 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n251), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n268), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n267), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n236), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n271), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n232) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_U31 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n250), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n276), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n271) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_U30 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n237), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n248), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n250) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_U29 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n239), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n272), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n236) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_U28 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n242), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n265), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n243), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n233) );
  AND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_U27 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n261), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n231), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n243) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_U26 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n276), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n248), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n265) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_U25 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n230), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n229), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n248) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_U24 ( .A(
        F_SD2_RedSB_inst_n73), .B(Red_StateRegOutput[99]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n230) );
  OR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_U23 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n261), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n231), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n242) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_U22 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n268), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n266), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n231) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_U21 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n228), .B(
        Red_StateRegOutput[98]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n268) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_U20 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n227), .B(
        F_SD2_RedSB_inst_n74), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n228) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_U19 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n267), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n270), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n261) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_U18 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n272), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n270) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_U17 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n226), .B(
        Red_StateRegOutput[101]), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n272) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_U16 ( .A(
        F_SD2_RedSB_inst_n73), .B(F_SD2_RedSB_inst_n76), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n226) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_U15 ( .A(
        Red_StateRegOutput[103]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n229), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n237) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_U14 ( .A(
        F_SD2_RedSB_inst_n76), .B(F_SD2_RedSB_inst_n74), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n229) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_U13 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n225), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n234) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_U12 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n267), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n239), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n224), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n225) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_U11 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n267), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n239), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n276), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n224) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_U10 ( .A(
        Red_StateRegOutput[100]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n227), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n276) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_U9 ( .A(
        F_SD2_RedSB_inst_n75), .B(F_SD2_RedSB_inst_n73), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n227) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_U8 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n266), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n239) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_U7 ( .A(
        Red_StateRegOutput[104]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n223), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n266) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_U6 ( .A(
        F_SD2_RedSB_inst_n75), .B(F_SD2_RedSB_inst_n76), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n223) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_U5 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n251), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n267) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_U4 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n222), .B(
        Red_StateRegOutput[102]), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n251) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_U3 ( .A(
        F_SD2_RedSB_inst_n75), .B(F_SD2_RedSB_inst_n74), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_104_n222) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_U69 ( .A(
        Red_StateRegOutput[106]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n280), .Z(Red_Feedback[0])
         );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_U68 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n279), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n278), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n280) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_U67 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n277), .B2(
        Red_StateRegOutput[107]), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n276), .C2(
        Red_StateRegOutput[110]), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n275), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n278) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_U66 ( .A1(
        Red_StateRegOutput[107]), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n277), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n276), .B2(
        Red_StateRegOutput[110]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n275) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_U65 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n274), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n273), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n276) );
  AOI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_U64 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n272), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n271), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n270), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n269), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n273) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_U63 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n268), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n267), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n266), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n265), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n264), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n269) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_U62 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n268), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n263), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n262), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n270) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_U61 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n268), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n263), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n261), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n262) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_U60 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n260), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n259), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n258), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n271) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_U59 ( .A(
        Red_StateRegOutput[105]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n257), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n274) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_U58 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n253), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n252), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n251), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n254) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_U57 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n252), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n253), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n250), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n255) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_U56 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n242), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n241), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n243), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n240), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n239), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n277) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_U55 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n238), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n237), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n236), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n239) );
  AOI222_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_U54 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n253), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n251), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n253), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n235), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n251), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n235), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n237) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_U53 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n245), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n267), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n235) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_U52 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n263), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n249), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n251) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_U51 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n234), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n253) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_U50 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n256), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n233), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n240) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_U49 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n261), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n263), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n232), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n241) );
  NOR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_U48 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n267), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n247), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n259), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n232) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_U47 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n248), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n249), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n259) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_U46 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n268), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n231), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n247) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_U45 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n256), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n267) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_U44 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n245), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n248), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n261) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_U43 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n264), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n260), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n230), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n279) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_U42 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n249), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n229), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n228), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n230) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_U41 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n249), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n227), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n250), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n228) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_U40 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n238), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n250) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_U39 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n245), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n265), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n238) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_U38 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n242), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n231), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n265) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_U37 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n244), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n246), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n256), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n263), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n227) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_U36 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n243), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n248), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n246) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_U35 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n266), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n245), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n244) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_U34 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n272), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n226), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n258), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n229) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_U33 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n234), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n225), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n258) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_U32 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n243), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n231), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n226) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_U31 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n234), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n225), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n260) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_U30 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n231), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n256), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n225) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_U29 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n224), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n223), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n256) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_U28 ( .A(
        Red_StateRegOutput[105]), .B(F_SD2_RedSB_inst_n77), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n224) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_U27 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n263), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n231) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_U26 ( .A(
        Red_StateRegOutput[111]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n222), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n263) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_U25 ( .A(
        F_SD2_RedSB_inst_n80), .B(F_SD2_RedSB_inst_n79), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n222) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_U24 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n242), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n268), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n234) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_U23 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n266), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n268) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_U22 ( .A(
        Red_StateRegOutput[109]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n223), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n266) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_U21 ( .A(
        F_SD2_RedSB_inst_n78), .B(F_SD2_RedSB_inst_n79), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n223) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_U20 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n243), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n242) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_U19 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n221), .B(
        Red_StateRegOutput[108]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n243) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_U18 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n233), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n264) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_U17 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n252), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n249), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n233) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_U16 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n220), .B(
        F_SD2_RedSB_inst_n78), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n249) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_U15 ( .A(
        Red_StateRegOutput[106]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n221), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n220) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_U14 ( .A(
        F_SD2_RedSB_inst_n80), .B(F_SD2_RedSB_inst_n77), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n221) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_U13 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n245), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n248), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n252) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_U12 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n236), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n248) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_U11 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n219), .B(
        Red_StateRegOutput[107]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n236) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_U10 ( .A(
        F_SD2_RedSB_inst_n77), .B(F_SD2_RedSB_inst_n79), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n219) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_U9 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n272), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n245) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_U8 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n218), .B(
        F_SD2_RedSB_inst_n78), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n272) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_U7 ( .A(
        Red_StateRegOutput[110]), .B(F_SD2_RedSB_inst_n80), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n218) );
  OAI33_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_U6 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n256), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n215), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n217), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n267), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n255), .B3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n254), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n257) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_U5 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n249), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n216), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n217) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_U4 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n245), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n246), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n243), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n244), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n216) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_U3 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n248), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n247), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_105_n215) );
  AOI222_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_U69 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n279), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n278), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n279), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n277), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n278), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n276), .ZN(Red_Feedback[1])
         );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_U68 ( .A(
        Red_StateRegOutput[110]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n275), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n276) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_U67 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n274), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n273), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n272), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n273), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n271), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n275) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_U66 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n270), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n269), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n268), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n269), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n267), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n271) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_U65 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n266), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n267) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_U64 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n265), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n264), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n268) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_U63 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n263), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n262), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n261), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n272) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_U62 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n260), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n259), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n262) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_U61 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n265), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n264), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n258), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n274) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_U60 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n265), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n264), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n257), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n258) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_U59 ( .A(
        Red_StateRegOutput[106]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n256), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n277) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_U58 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n255), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n254), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n253), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n256) );
  AOI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_U57 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n266), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n252), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n251), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n250), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n253) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_U56 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n249), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n248), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n260), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n261), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n250) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_U55 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n247), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n246), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n261) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_U54 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n245), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n260), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n244), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n243), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n249) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_U53 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n242), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n260) );
  NOR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_U52 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n241), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n240), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n239), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n251) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_U51 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n263), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n252) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_U50 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n247), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n246), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n263) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_U49 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n265), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n238), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n246) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_U48 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n244), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n238), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n254) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_U47 ( .A(
        Red_StateRegOutput[105]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n237), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n278) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_U46 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n238), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n236), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n235), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n237) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_U45 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n238), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n234), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n233), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n235) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_U44 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n244), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n247), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n259), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n248), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n233) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_U43 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n232), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n264), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n239), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n255), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n236) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_U42 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n257), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n241), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n255) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_U41 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n257), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n265), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n242), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n231), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n232) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_U40 ( .A(
        Red_StateRegOutput[107]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n230), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n279) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_U39 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n229), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n259), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n228), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n257), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n227), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n230) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_U38 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n226), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n225), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n224), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n223), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n227) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_U37 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n257), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n244), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n223) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_U36 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n222), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n224) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_U35 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n241), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n266), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n225) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_U34 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n257), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n239), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n266) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_U33 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n242), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n248), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n239) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_U32 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n259), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n257) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_U31 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n234), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n221), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n228) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_U30 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n222), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n247), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n231), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n240), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n221) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_U29 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n241), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n248), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n231) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_U28 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n273), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n248) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_U27 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n273), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n238), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n222) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_U26 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n273), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n245), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n244), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n247), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n234) );
  AND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_U25 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n270), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n264), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n247) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_U24 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n265), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n242), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n244) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_U23 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n240), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n265) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_U22 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n240), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n270), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n245) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_U21 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n241), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n270) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_U20 ( .A(
        Red_StateRegOutput[110]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n220), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n273) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_U19 ( .A(
        F_SD2_RedSB_inst_n79), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n219), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n259) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_U18 ( .A(
        Red_StateRegOutput[107]), .B(F_SD2_RedSB_inst_n77), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n219) );
  NOR4_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_U17 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n242), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n241), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n240), .A4(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n269), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n229) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_U16 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n243), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n269) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_U15 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n264), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n226), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n243) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_U14 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n238), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n226) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_U13 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n218), .B(
        Red_StateRegOutput[105]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n238) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_U12 ( .A(
        F_SD2_RedSB_inst_n77), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n217), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n218) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_U11 ( .A(
        Red_StateRegOutput[109]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n217), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n264) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_U10 ( .A(
        F_SD2_RedSB_inst_n79), .B(F_SD2_RedSB_inst_n78), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n217) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_U9 ( .A(
        Red_StateRegOutput[111]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n216), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n240) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_U8 ( .A(
        F_SD2_RedSB_inst_n79), .B(F_SD2_RedSB_inst_n80), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n216) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_U7 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n215), .B(
        Red_StateRegOutput[108]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n241) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_U6 ( .A(
        F_SD2_RedSB_inst_n77), .B(F_SD2_RedSB_inst_n80), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n215) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_U5 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n214), .B(
        Red_StateRegOutput[106]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n242) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_U4 ( .A(
        F_SD2_RedSB_inst_n77), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n220), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n214) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_U3 ( .A(
        F_SD2_RedSB_inst_n78), .B(F_SD2_RedSB_inst_n80), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_106_n220) );
  MUX2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_U54 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n240), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n239), .S(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n238), .Z(Red_Feedback[2])
         );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_U53 ( .A(
        Red_StateRegOutput[107]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n237), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n238) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_U52 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n236), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n235), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n234), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n233), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n237) );
  OR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_U51 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n232), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n231), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n230), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n233) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_U50 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n229), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n228), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n227), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n234) );
  AOI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_U49 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n226), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n225), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n224), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n223), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n236) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_U48 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n222), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n221), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n220), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n221), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n219), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n223) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_U47 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n226), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n225), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n218), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n221) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_U46 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n217), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n216), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n225) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_U45 ( .A(
        Red_StateRegOutput[110]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n215), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n239) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_U44 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n214), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n230), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n213), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n212), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n215) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_U43 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n228), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n226), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n211), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n232), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n212) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_U42 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n210), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n228), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n210), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n226), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n216), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n213) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_U41 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n220), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n216) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_U40 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n209), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n226) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_U39 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n208), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n207), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n228) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_U38 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n219), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n206), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n205), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n210) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_U37 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n219), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n206), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n208), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n205) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_U36 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n235), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n208) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_U35 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n222), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n204), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n229), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n214) );
  AND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_U34 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n206), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n219), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n204) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_U33 ( .A(
        Red_StateRegOutput[106]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n203), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n240) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_U32 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n202), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n201), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n200), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n201), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n199), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n203) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_U31 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n198), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n197), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n230), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n209), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n199) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_U30 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n227), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n220), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n218), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n197) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_U29 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n207), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n218) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_U28 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n222), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n201), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n227) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_U27 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n198), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n230), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n209), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n230), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n217), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n200) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_U26 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n231), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n206), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n209) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_U25 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n207), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n235), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n220), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n230) );
  AOI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_U24 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n229), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n211), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n207), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n224), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n198) );
  NOR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_U23 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n231), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n220), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n201), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n224) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_U22 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n219), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n220), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n211) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_U21 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n196), .B(
        Red_StateRegOutput[110]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n220) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_U20 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n201), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n219) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_U19 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n232), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n206), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n229) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_U18 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n195), .B(
        Red_StateRegOutput[109]), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n206) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_U17 ( .A(
        F_SD2_RedSB_inst_n79), .B(F_SD2_RedSB_inst_n78), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n195) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_U16 ( .A(
        Red_StateRegOutput[111]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n194), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n201) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_U15 ( .A(
        F_SD2_RedSB_inst_n79), .B(F_SD2_RedSB_inst_n80), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n194) );
  NOR4_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_U14 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n207), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n231), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n232), .A4(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n235), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n202) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_U13 ( .A(
        Red_StateRegOutput[107]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n193), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n235) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_U12 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n217), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n232) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_U11 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n192), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n193), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n217) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_U10 ( .A(
        F_SD2_RedSB_inst_n77), .B(F_SD2_RedSB_inst_n79), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n193) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_U9 ( .A(
        F_SD2_RedSB_inst_n78), .B(Red_StateRegOutput[105]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n192) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_U8 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n222), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n231) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_U7 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n191), .B(
        Red_StateRegOutput[108]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n222) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_U6 ( .A(
        F_SD2_RedSB_inst_n77), .B(F_SD2_RedSB_inst_n80), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n191) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_U5 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n190), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n196), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n207) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_U4 ( .A(
        F_SD2_RedSB_inst_n78), .B(F_SD2_RedSB_inst_n80), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n196) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_U3 ( .A(
        F_SD2_RedSB_inst_n77), .B(Red_StateRegOutput[106]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_107_n190) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_U70 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n290), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n289), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n288), .ZN(Red_Feedback[3])
         );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_U69 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n290), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n287), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n288) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_U68 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n286), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n285), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n284), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n287) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_U67 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n283), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n282), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n286), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n284) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_U66 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n289), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n285) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_U65 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n283), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n282), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n281), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n289) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_U64 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n282), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n286), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n283), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n281) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_U63 ( .A(
        Red_StateRegOutput[110]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n268), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n282) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_U62 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n267), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n266), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n265), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n269), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n268) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_U61 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n264), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n274), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n263), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n262), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n261), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n265) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_U60 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n260), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n259), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n278), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n258), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n263) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_U59 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n262), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n274) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_U58 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n273), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n272), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n264) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_U57 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n257), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n266) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_U56 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n256), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n255), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n254), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n267) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_U55 ( .A(
        Red_StateRegOutput[107]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n253), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n283) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_U54 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n252), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n262), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n251), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n250), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n253) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_U53 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n278), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n257), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n249), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n250) );
  NAND4_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_U52 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n254), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n248), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n276), .A4(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n262), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n251) );
  AOI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_U51 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n271), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n247), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n246), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n277), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n252) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_U50 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n258), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n259), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n245), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n277) );
  NOR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_U49 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n278), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n244), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n280), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n246) );
  AND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_U48 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n258), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n259), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n280) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_U47 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n243), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n259) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_U46 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n249), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n269), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n271) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_U45 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n242), .B(
        Red_StateRegOutput[106]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n290) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_U44 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n276), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n279), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n257) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_U43 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n262), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n269), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n279) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_U42 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n244), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n256), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n245) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_U41 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n240), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n247), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n256) );
  AND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_U40 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n243), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n241), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n261) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_U39 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n278), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n272), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n241) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_U38 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n249), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n273), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n243) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_U37 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n255), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n273) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_U36 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n249), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n247), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n248) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_U35 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n275), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n255), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n254) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_U34 ( .A(
        Red_StateRegOutput[109]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n239), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n255) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_U33 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n278), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n275) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_U32 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n269), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n244) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_U31 ( .A(
        Red_StateRegOutput[110]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n238), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n269) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_U30 ( .A(
        F_SD2_RedSB_inst_n78), .B(F_SD2_RedSB_inst_n80), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n238) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_U29 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n262), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n240), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n270) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_U28 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n249), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n240) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_U27 ( .A(
        Red_StateRegOutput[108]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n237), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n249) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_U26 ( .A(
        F_SD2_RedSB_inst_n77), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n236), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n262) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_U25 ( .A(
        Red_StateRegOutput[107]), .B(F_SD2_RedSB_inst_n79), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n236) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_U24 ( .A(
        F_SD2_RedSB_inst_n78), .B(F_SD2_RedSB_inst_n79), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n239) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_U23 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n276), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n247), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n258) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_U22 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n272), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n247) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_U21 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n235), .B(
        Red_StateRegOutput[111]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n272) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_U20 ( .A(
        F_SD2_RedSB_inst_n79), .B(F_SD2_RedSB_inst_n80), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n235) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_U19 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n260), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n276) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_U18 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n234), .B(
        Red_StateRegOutput[106]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n260) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_U17 ( .A(
        F_SD2_RedSB_inst_n78), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n237), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n234) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_U16 ( .A(
        F_SD2_RedSB_inst_n77), .B(F_SD2_RedSB_inst_n80), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n237) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_U15 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n258), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n230), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n232), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n233), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n242) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_U14 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n261), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n269), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n261), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n248), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n260), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n233) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_U13 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n243), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n257), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n241), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n257), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n231), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n232) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_U12 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n260), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n245), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n231) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_U11 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n278), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n270), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n244), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n254), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n230) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_U10 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n229), .B(
        Red_StateRegOutput[105]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n286) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_U9 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n225), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n277), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n228), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n229) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_U8 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n276), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n226), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n275), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n227), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n228) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_U7 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n274), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n272), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n273), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n227) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_U6 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n269), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n270), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n273), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n271), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n226) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_U5 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n280), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n279), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n278), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n225) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_U4 ( .A(
        Red_StateRegOutput[105]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n224), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n278) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_U3 ( .A(
        F_SD2_RedSB_inst_n77), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n239), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_108_n224) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_U73 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n282), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n281), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n282), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n280), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n279), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n283) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_U72 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n278), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n277), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n276), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n284) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_U71 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n275), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n274), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n277), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n276) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_U70 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n273), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n272), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n271), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n275) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_U69 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n270), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n277) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_U68 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n264), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n263), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n262), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n265) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_U67 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n263), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n267) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_U66 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n278), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n261) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_U65 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n259), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n258), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n278) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_U64 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n262), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n279), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n256), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n274) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_U63 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n281), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n273), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n257) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_U62 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n262), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n255), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n281) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_U61 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n272), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n280), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n263), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n252), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n253) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_U60 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n259), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n260), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n251), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n285), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n252) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_U59 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n270), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n250), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n285) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_U58 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n268), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n249), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n280) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_U57 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n286), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n272) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_U56 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n255), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n248), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n286) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_U55 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n247), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n246), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n245), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n254) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_U54 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n258), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n269), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n247), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n245) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_U53 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n271), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n244), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n243), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n246) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_U52 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n282), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n243) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_U51 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n268), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n249), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n282) );
  OR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_U50 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n273), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n250), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n249) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_U49 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n264), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n268) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_U48 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n251), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n273), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n244) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_U47 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n279), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n251) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_U46 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n270), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n241), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n240), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n242) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_U45 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n258), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n260), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n239), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n238), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n240) );
  OR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_U44 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n247), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n269), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n266), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n238) );
  OR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_U43 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n279), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n250), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n259), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n266) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_U42 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n255), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n247) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_U41 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n264), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n248), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n263), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n237), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n250), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n239) );
  AND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_U40 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n264), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n248), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n237) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_U39 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n273), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n255), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n263) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_U38 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n262), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n279), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n248) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_U37 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n259), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n262) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_U36 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n270), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n271), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n264) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_U35 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n271), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n250), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n260) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_U34 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n269), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n271) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_U33 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n273), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n279), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n258) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_U32 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n256), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n273) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_U31 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n256), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n236), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n259), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n236), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n250), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n241) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_U30 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n235), .B(
        Red_StateRegOutput[105]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n250) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_U29 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n234), .B(
        F_SD2_RedSB_inst_n78), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n235) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_U28 ( .A(
        Red_StateRegOutput[107]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n234), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n259) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_U27 ( .A(
        F_SD2_RedSB_inst_n79), .B(F_SD2_RedSB_inst_n77), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n234) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_U26 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n255), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n279), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n269), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n236) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_U25 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n233), .B(
        Red_StateRegOutput[108]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n269) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_U24 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n232), .B(
        F_SD2_RedSB_inst_n78), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n279) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_U23 ( .A(
        Red_StateRegOutput[110]), .B(F_SD2_RedSB_inst_n80), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n232) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_U22 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n231), .B(
        Red_StateRegOutput[106]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n255) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_U21 ( .A(
        F_SD2_RedSB_inst_n78), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n233), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n231) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_U20 ( .A(
        F_SD2_RedSB_inst_n77), .B(F_SD2_RedSB_inst_n80), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n233) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_U19 ( .A(
        Red_StateRegOutput[111]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n230), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n256) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_U18 ( .A(
        F_SD2_RedSB_inst_n79), .B(F_SD2_RedSB_inst_n80), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n230) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_U17 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n229), .B(
        Red_StateRegOutput[109]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n270) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_U16 ( .A(
        F_SD2_RedSB_inst_n79), .B(F_SD2_RedSB_inst_n78), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n229) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_U15 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n217), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n219), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n227), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n221), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n228), .ZN(Red_Feedback[4])
         );
  NOR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_U14 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n219), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n221), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n227), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n228) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_U13 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n225), .B2(
        Red_StateRegOutput[107]), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n226), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n227) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_U12 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n225), .B2(
        Red_StateRegOutput[107]), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n217), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n226) );
  AOI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_U11 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n269), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n222), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n223), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n224), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n225) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_U10 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n286), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n260), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n261), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n269), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n224) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_U9 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n265), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n266), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n267), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n268), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n223) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_U8 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n285), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n257), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n274), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n222) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_U7 ( .A(
        Red_StateRegOutput[110]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n220), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n221) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_U6 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n286), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n285), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n284), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n283), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n220) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_U5 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n218), .B(
        Red_StateRegOutput[106]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n219) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_U4 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n254), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n253), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n218) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_U3 ( .A(
        Red_StateRegOutput[105]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n242), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_109_n217) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_U72 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n283), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n282), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n281), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n280), .ZN(Red_Feedback[5])
         );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_U71 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n279), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n280), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n278), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n282) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_U70 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n279), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n280), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n281), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n278) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_U69 ( .A(
        Red_StateRegOutput[110]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n277), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n281) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_U68 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n276), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n275), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n277) );
  NAND4_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_U67 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n274), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n273), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n272), .A4(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n271), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n275) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_U66 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n270), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n269), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n268), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n267), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n276) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_U65 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n266), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n267) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_U64 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n273), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n265), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n264), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n263), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n269) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_U63 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n262), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n264) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_U62 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n261), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n271), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n260), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n259), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n265) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_U61 ( .A(
        Red_StateRegOutput[106]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n258), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n280) );
  NOR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_U60 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n257), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n256), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n255), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n258) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_U59 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n253), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n252), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n262) );
  AOI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_U58 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n274), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n251), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n250), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n249), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n256) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_U57 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n248), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n247), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n274), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n249) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_U56 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n270), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n246), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n251) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_U55 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n247), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n270) );
  NOR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_U54 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n253), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n246), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n252), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n257) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_U53 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n259), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n250), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n252) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_U52 ( .A(
        Red_StateRegOutput[105]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n245), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n279) );
  AOI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_U51 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n274), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n244), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n243), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n242), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n245) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_U50 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n253), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n241), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n254), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n240), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n242) );
  OR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_U49 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n253), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n241), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n259), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n240) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_U48 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n239), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n250), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n246), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n254) );
  NOR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_U47 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n239), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n238), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n271), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n243) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_U46 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n273), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n261), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n248), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n237), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n238) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_U45 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n236), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n259), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n235), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n244) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_U44 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n234), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n248), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n261), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n235) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_U43 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n233), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n236) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_U42 ( .A(
        Red_StateRegOutput[107]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n232), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n283) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_U41 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n261), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n231), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n230), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n232) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_U40 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n266), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n229), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n228), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n263), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n230) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_U39 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n246), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n227), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n263) );
  NAND4_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_U38 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n239), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n268), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n273), .A4(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n229), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n228) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_U37 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n271), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n268) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_U36 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n239), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n272), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n261), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n233), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n266) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_U35 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n247), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n250), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n233) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_U34 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n246), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n241), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n272) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_U33 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n247), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n227), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n241) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_U32 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n259), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n239) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_U31 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n273), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n226), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n225), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n253), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n231) );
  AOI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_U30 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n234), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n246), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n260), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n246), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n237), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n226) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_U29 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n274), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n247), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n237) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_U28 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n229), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n274) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_U27 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n253), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n260) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_U26 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n229), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n271), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n253) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_U25 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n224), .B(
        Red_StateRegOutput[109]), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n271) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_U24 ( .A(
        F_SD2_RedSB_inst_n78), .B(F_SD2_RedSB_inst_n79), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n224) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_U23 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n223), .B(
        Red_StateRegOutput[108]), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n229) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_U22 ( .A(
        F_SD2_RedSB_inst_n77), .B(F_SD2_RedSB_inst_n80), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n223) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_U21 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n248), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n246) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_U20 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n222), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n221), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n248) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_U19 ( .A(
        F_SD2_RedSB_inst_n80), .B(Red_StateRegOutput[106]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n222) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_U18 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n225), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n234) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_U17 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n259), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n247), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n225) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_U16 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n220), .B(
        Red_StateRegOutput[110]), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n247) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_U15 ( .A(
        F_SD2_RedSB_inst_n78), .B(F_SD2_RedSB_inst_n80), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n220) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_U14 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n219), .B(
        F_SD2_RedSB_inst_n79), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n259) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_U13 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n221), .B(
        Red_StateRegOutput[105]), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n219) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_U12 ( .A(
        F_SD2_RedSB_inst_n77), .B(F_SD2_RedSB_inst_n78), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n221) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_U11 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n250), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n273) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_U10 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n218), .B(
        Red_StateRegOutput[111]), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n250) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_U9 ( .A(
        F_SD2_RedSB_inst_n79), .B(F_SD2_RedSB_inst_n80), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n218) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_U8 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n227), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n261) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_U7 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n217), .B(
        F_SD2_RedSB_inst_n79), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n227) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_U6 ( .A(
        Red_StateRegOutput[107]), .B(F_SD2_RedSB_inst_n77), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n217) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_U5 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n254), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n215), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n216), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n255) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_U4 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n272), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n262), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n216) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_U3 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n268), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n270), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n261), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n274), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_110_n215) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_U65 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n283), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n282), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n281), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n280), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n279), .ZN(Red_Feedback[6])
         );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_U64 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n283), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n282), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n281), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n279) );
  MUX2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_U63 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n283), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n282), .S(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n278), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n280) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_U62 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n277), .B(
        Red_StateRegOutput[107]), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n278) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_U61 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n276), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n275), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n274), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n277) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_U60 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n273), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n274) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_U59 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n272), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n271), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n270), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n269), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n268), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n273) );
  AND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_U58 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n267), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n266), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n265), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n269) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_U57 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n266), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n264), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n263), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n262), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n275) );
  AOI222_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_U56 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n261), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n260), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n261), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n259), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n260), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n259), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n263) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_U55 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n258), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n268), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n259) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_U54 ( .A(
        Red_StateRegOutput[105]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n257), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n281) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_U53 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n268), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n256), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n255), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n257) );
  NAND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_U52 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n268), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n254), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n262), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n255) );
  AOI222_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_U51 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n261), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n260), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n261), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n253), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n260), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n253), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n254) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_U50 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n276), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n258), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n253) );
  OAI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_U49 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n252), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n251), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n250), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n249), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n256) );
  AOI22_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_U48 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n276), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n266), .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n248), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n247), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n252) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_U47 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n264), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n247) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_U46 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n272), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n258), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n264) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_U45 ( .A(
        Red_StateRegOutput[106]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n246), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n282) );
  OAI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_U44 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n248), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n262), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n245), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n244), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n246) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_U43 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n248), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n243), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n244) );
  AOI211_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_U42 ( .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n271), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n242), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n241), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n240), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n245) );
  NOR3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_U41 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n270), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n239), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n250), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n240) );
  AND3_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_U40 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n238), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n268), .A3(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n260), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n241) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_U39 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n248), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n266), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n260) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_U38 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n251), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n237), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n249), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n238) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_U37 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n276), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n270), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n249) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_U36 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n258), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n236), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n262) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_U35 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n237), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n258) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_U34 ( .A(
        Red_StateRegOutput[110]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n235), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n283) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_U33 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n234), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n237), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n233), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n237), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n232), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n235) );
  OAI221_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_U32 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n251), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n268), .C1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n267), .C2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n236), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n271), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n232) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_U31 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n250), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n276), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n271) );
  NAND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_U30 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n237), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n248), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n250) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_U29 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n239), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n272), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n236) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_U28 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n242), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n265), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n243), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n233) );
  AND2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_U27 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n261), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n231), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n243) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_U26 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n276), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n248), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n265) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_U25 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n230), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n229), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n248) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_U24 ( .A(
        F_SD2_RedSB_inst_n77), .B(Red_StateRegOutput[106]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n230) );
  OR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_U23 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n261), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n231), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n242) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_U22 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n268), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n266), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n231) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_U21 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n228), .B(
        Red_StateRegOutput[105]), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n268) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_U20 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n227), .B(
        F_SD2_RedSB_inst_n78), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n228) );
  NOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_U19 ( .A1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n267), .A2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n270), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n261) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_U18 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n272), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n270) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_U17 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n226), .B(
        Red_StateRegOutput[108]), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n272) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_U16 ( .A(
        F_SD2_RedSB_inst_n77), .B(F_SD2_RedSB_inst_n80), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n226) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_U15 ( .A(
        Red_StateRegOutput[110]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n229), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n237) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_U14 ( .A(
        F_SD2_RedSB_inst_n80), .B(F_SD2_RedSB_inst_n78), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n229) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_U13 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n225), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n234) );
  AOI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_U12 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n267), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n239), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n224), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n225) );
  OAI21_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_U11 ( .B1(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n267), .B2(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n239), .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n276), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n224) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_U10 ( .A(
        Red_StateRegOutput[107]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n227), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n276) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_U9 ( .A(
        F_SD2_RedSB_inst_n79), .B(F_SD2_RedSB_inst_n77), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n227) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_U8 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n266), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n239) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_U7 ( .A(
        Red_StateRegOutput[111]), .B(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n223), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n266) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_U6 ( .A(
        F_SD2_RedSB_inst_n79), .B(F_SD2_RedSB_inst_n80), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n223) );
  INV_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_U5 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n251), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n267) );
  XOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_U4 ( .A(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n222), .B(
        Red_StateRegOutput[109]), .Z(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n251) );
  XNOR2_X1 F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_U3 ( .A(
        F_SD2_RedSB_inst_n79), .B(F_SD2_RedSB_inst_n78), .ZN(
        F_SD2_RedSB_inst_F_SD2_RedSB_bit_inst_111_n222) );
  BUF_X1 K0K1_KeyMUX_And_Red_KeyMUX_U32 ( .A(n3), .Z(
        K0K1_KeyMUX_And_Red_KeyMUX_n67) );
  BUF_X1 K0K1_KeyMUX_And_Red_KeyMUX_U31 ( .A(n4), .Z(
        K0K1_KeyMUX_And_Red_KeyMUX_n74) );
  BUF_X2 K0K1_KeyMUX_And_Red_KeyMUX_U30 ( .A(n7), .Z(
        K0K1_KeyMUX_And_Red_KeyMUX_n89) );
  BUF_X1 K0K1_KeyMUX_And_Red_KeyMUX_U29 ( .A(n3), .Z(
        K0K1_KeyMUX_And_Red_KeyMUX_n66) );
  BUF_X1 K0K1_KeyMUX_And_Red_KeyMUX_U28 ( .A(n3), .Z(
        K0K1_KeyMUX_And_Red_KeyMUX_n65) );
  BUF_X1 K0K1_KeyMUX_And_Red_KeyMUX_U27 ( .A(n4), .Z(
        K0K1_KeyMUX_And_Red_KeyMUX_n73) );
  BUF_X1 K0K1_KeyMUX_And_Red_KeyMUX_U26 ( .A(n3), .Z(
        K0K1_KeyMUX_And_Red_KeyMUX_n68) );
  BUF_X4 K0K1_KeyMUX_And_Red_KeyMUX_U25 ( .A(K0K1_KeyMUX_And_Red_KeyMUX_n65), 
        .Z(K0K1_KeyMUX_And_Red_KeyMUX_n69) );
  BUF_X2 K0K1_KeyMUX_And_Red_KeyMUX_U24 ( .A(n4), .Z(
        K0K1_KeyMUX_And_Red_KeyMUX_n82) );
  BUF_X2 K0K1_KeyMUX_And_Red_KeyMUX_U23 ( .A(K0K1_KeyMUX_And_Red_KeyMUX_n89), 
        .Z(K0K1_KeyMUX_And_Red_KeyMUX_n88) );
  BUF_X4 K0K1_KeyMUX_And_Red_KeyMUX_U22 ( .A(K0K1_KeyMUX_And_Red_KeyMUX_n88), 
        .Z(K0K1_KeyMUX_And_Red_KeyMUX_n86) );
  CLKBUF_X3 K0K1_KeyMUX_And_Red_KeyMUX_U21 ( .A(n5), .Z(
        K0K1_KeyMUX_And_Red_KeyMUX_n58) );
  BUF_X8 K0K1_KeyMUX_And_Red_KeyMUX_U20 ( .A(K0K1_KeyMUX_And_Red_KeyMUX_n58), 
        .Z(K0K1_KeyMUX_And_Red_KeyMUX_n62) );
  BUF_X4 K0K1_KeyMUX_And_Red_KeyMUX_U19 ( .A(K0K1_KeyMUX_And_Red_KeyMUX_n59), 
        .Z(K0K1_KeyMUX_And_Red_KeyMUX_n61) );
  BUF_X2 K0K1_KeyMUX_And_Red_KeyMUX_U18 ( .A(K0K1_KeyMUX_And_Red_KeyMUX_n89), 
        .Z(K0K1_KeyMUX_And_Red_KeyMUX_n85) );
  BUF_X4 K0K1_KeyMUX_And_Red_KeyMUX_U17 ( .A(K0K1_KeyMUX_And_Red_KeyMUX_n85), 
        .Z(K0K1_KeyMUX_And_Red_KeyMUX_n87) );
  CLKBUF_X3 K0K1_KeyMUX_And_Red_KeyMUX_U16 ( .A(K0K1_KeyMUX_And_Red_KeyMUX_n59), .Z(K0K1_KeyMUX_And_Red_KeyMUX_n60) );
  CLKBUF_X3 K0K1_KeyMUX_And_Red_KeyMUX_U15 ( .A(K0K1_KeyMUX_And_Red_KeyMUX_n58), .Z(K0K1_KeyMUX_And_Red_KeyMUX_n63) );
  BUF_X4 K0K1_KeyMUX_And_Red_KeyMUX_U14 ( .A(K0K1_KeyMUX_And_Red_KeyMUX_n67), 
        .Z(K0K1_KeyMUX_And_Red_KeyMUX_n71) );
  BUF_X4 K0K1_KeyMUX_And_Red_KeyMUX_U13 ( .A(K0K1_KeyMUX_And_Red_KeyMUX_n66), 
        .Z(K0K1_KeyMUX_And_Red_KeyMUX_n70) );
  BUF_X2 K0K1_KeyMUX_And_Red_KeyMUX_U12 ( .A(n7), .Z(
        K0K1_KeyMUX_And_Red_KeyMUX_n83) );
  CLKBUF_X3 K0K1_KeyMUX_And_Red_KeyMUX_U11 ( .A(K0K1_KeyMUX_And_Red_KeyMUX_n68), .Z(K0K1_KeyMUX_And_Red_KeyMUX_n72) );
  BUF_X2 K0K1_KeyMUX_And_Red_KeyMUX_U10 ( .A(K0K1_KeyMUX_And_Red_KeyMUX_n74), 
        .Z(K0K1_KeyMUX_And_Red_KeyMUX_n75) );
  BUF_X2 K0K1_KeyMUX_And_Red_KeyMUX_U9 ( .A(K0K1_KeyMUX_And_Red_KeyMUX_n73), 
        .Z(K0K1_KeyMUX_And_Red_KeyMUX_n76) );
  BUF_X2 K0K1_KeyMUX_And_Red_KeyMUX_U8 ( .A(K0K1_KeyMUX_And_Red_KeyMUX_n89), 
        .Z(K0K1_KeyMUX_And_Red_KeyMUX_n84) );
  BUF_X2 K0K1_KeyMUX_And_Red_KeyMUX_U7 ( .A(K0K1_KeyMUX_And_Red_KeyMUX_n73), 
        .Z(K0K1_KeyMUX_And_Red_KeyMUX_n79) );
  BUF_X2 K0K1_KeyMUX_And_Red_KeyMUX_U6 ( .A(K0K1_KeyMUX_And_Red_KeyMUX_n74), 
        .Z(K0K1_KeyMUX_And_Red_KeyMUX_n80) );
  BUF_X2 K0K1_KeyMUX_And_Red_KeyMUX_U5 ( .A(K0K1_KeyMUX_And_Red_KeyMUX_n74), 
        .Z(K0K1_KeyMUX_And_Red_KeyMUX_n77) );
  BUF_X2 K0K1_KeyMUX_And_Red_KeyMUX_U4 ( .A(K0K1_KeyMUX_And_Red_KeyMUX_n73), 
        .Z(K0K1_KeyMUX_And_Red_KeyMUX_n78) );
  BUF_X32 K0K1_KeyMUX_And_Red_KeyMUX_U3 ( .A(n6), .Z(
        K0K1_KeyMUX_And_Red_KeyMUX_n64) );
  BUF_X2 K0K1_KeyMUX_And_Red_KeyMUX_U2 ( .A(K0K1_KeyMUX_And_Red_KeyMUX_n73), 
        .Z(K0K1_KeyMUX_And_Red_KeyMUX_n81) );
  BUF_X4 K0K1_KeyMUX_And_Red_KeyMUX_U1 ( .A(n5), .Z(
        K0K1_KeyMUX_And_Red_KeyMUX_n59) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_0_U9 ( .A(KeyMux_D0_input[0]), 
        .B(KeyMux_D1_input[0]), .S(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_0_n30), .Z(Red_SelectedKey[0])
         );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_0_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_0_n29), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_0_n28), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_0_n27), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_0_n30) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_0_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n74), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_0_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n85), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_0_n27) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_0_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n74), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_0_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n85), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_0_n28) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_0_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_0_n25), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n68), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_0_n26) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_0_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_0_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_0_n25) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_0_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n68), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_0_n23), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_0_n29) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_0_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_0_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_0_n23) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_0_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_0_n24) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_1_U9 ( .A(KeyMux_D0_input[1]), 
        .B(KeyMux_D1_input[1]), .S(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_1_n30), .Z(Red_SelectedKey[1])
         );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_1_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_1_n29), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_1_n28), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_1_n27), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_1_n30) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_1_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n79), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_1_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n83), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_1_n27) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_1_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n79), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_1_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n83), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_1_n28) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_1_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_1_n25), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n68), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_1_n26) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_1_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_1_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_1_n25) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_1_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n68), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_1_n23), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_1_n29) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_1_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_1_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_1_n23) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_1_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_1_n24) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_2_U9 ( .A(KeyMux_D0_input[2]), 
        .B(KeyMux_D1_input[2]), .S(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_2_n30), .Z(Red_SelectedKey[2])
         );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_2_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_2_n29), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_2_n28), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_2_n27), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_2_n30) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_2_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n75), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_2_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n83), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_2_n27) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_2_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n75), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_2_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n83), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_2_n28) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_2_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_2_n25), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n69), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_2_n26) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_2_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n58), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_2_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_2_n25) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_2_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n69), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_2_n23), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n58), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_2_n29) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_2_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_2_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_2_n23) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_2_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n58), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_2_n24) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_3_U9 ( .A(KeyMux_D0_input[3]), 
        .B(KeyMux_D1_input[3]), .S(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_3_n31), .Z(Red_SelectedKey[3])
         );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_3_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_3_n30), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_3_n29), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_3_n28), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_3_n31) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_3_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n75), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_3_n27), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n83), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_3_n28) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_3_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n75), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_3_n27), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n83), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_3_n29) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_3_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_3_n26), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n69), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_3_n27) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_3_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n59), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_3_n25), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_3_n26) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_3_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n69), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_3_n24), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n59), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_3_n30) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_3_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_3_n25), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_3_n24) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_3_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n59), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_3_n25) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_4_U9 ( .A(KeyMux_D0_input[4]), 
        .B(KeyMux_D1_input[4]), .S(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_4_n31), .Z(Red_SelectedKey[4])
         );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_4_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_4_n30), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_4_n29), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_4_n28), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_4_n31) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_4_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n75), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_4_n27), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n83), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_4_n28) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_4_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n75), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_4_n27), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n83), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_4_n29) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_4_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_4_n26), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n69), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_4_n27) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_4_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n59), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_4_n25), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_4_n26) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_4_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n69), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_4_n24), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n59), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_4_n30) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_4_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_4_n25), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_4_n24) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_4_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n59), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_4_n25) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_5_U9 ( .A(KeyMux_D0_input[5]), 
        .B(KeyMux_D1_input[5]), .S(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_5_n30), .Z(Red_SelectedKey[5])
         );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_5_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_5_n29), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_5_n28), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_5_n27), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_5_n30) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_5_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n75), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_5_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n83), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_5_n27) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_5_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n75), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_5_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n83), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_5_n28) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_5_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_5_n25), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n69), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_5_n26) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_5_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n58), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_5_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_5_n25) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_5_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n69), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_5_n23), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n58), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_5_n29) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_5_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_5_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_5_n23) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_5_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n58), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_5_n24) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_6_U9 ( .A(KeyMux_D0_input[6]), 
        .B(KeyMux_D1_input[6]), .S(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_6_n30), .Z(Red_SelectedKey[6])
         );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_6_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_6_n29), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_6_n28), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_6_n27), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_6_n30) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_6_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n75), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_6_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n83), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_6_n27) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_6_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n75), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_6_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n83), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_6_n28) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_6_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_6_n25), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n69), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_6_n26) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_6_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n58), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_6_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_6_n25) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_6_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n69), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_6_n23), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n58), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_6_n29) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_6_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_6_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_6_n23) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_6_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n58), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_6_n24) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_7_U9 ( .A(KeyMux_D0_input[7]), 
        .B(KeyMux_D1_input[7]), .S(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_7_n31), .Z(Red_SelectedKey[7])
         );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_7_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_7_n30), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_7_n29), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_7_n28), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_7_n31) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_7_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n75), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_7_n27), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n83), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_7_n28) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_7_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n75), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_7_n27), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n83), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_7_n29) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_7_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_7_n26), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n69), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_7_n27) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_7_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n59), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_7_n25), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_7_n26) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_7_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n69), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_7_n24), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n59), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_7_n30) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_7_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_7_n25), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_7_n24) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_7_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n59), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_7_n25) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_8_U9 ( .A(KeyMux_D0_input[8]), 
        .B(KeyMux_D1_input[8]), .S(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_8_n31), .Z(Red_SelectedKey[8])
         );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_8_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_8_n30), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_8_n29), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_8_n28), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_8_n31) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_8_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n75), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_8_n27), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n83), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_8_n28) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_8_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n75), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_8_n27), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n83), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_8_n29) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_8_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_8_n26), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n69), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_8_n27) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_8_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n59), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_8_n25), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_8_n26) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_8_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n69), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_8_n24), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n59), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_8_n30) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_8_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_8_n25), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_8_n24) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_8_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n59), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_8_n25) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_9_U9 ( .A(KeyMux_D0_input[9]), 
        .B(KeyMux_D1_input[9]), .S(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_9_n30), .Z(Red_SelectedKey[9])
         );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_9_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_9_n29), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_9_n28), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_9_n27), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_9_n30) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_9_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n75), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_9_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n83), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_9_n27) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_9_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n75), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_9_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n83), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_9_n28) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_9_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_9_n25), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n69), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_9_n26) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_9_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n58), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_9_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_9_n25) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_9_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n69), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_9_n23), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n58), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_9_n29) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_9_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_9_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_9_n23) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_9_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n58), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_9_n24) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_10_U9 ( .A(
        KeyMux_D0_input[10]), .B(KeyMux_D1_input[10]), .S(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_10_n31), .Z(Red_SelectedKey[10]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_10_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_10_n30), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_10_n29), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_10_n28), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_10_n31) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_10_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n75), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_10_n27), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n83), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_10_n28) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_10_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n75), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_10_n27), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n83), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_10_n29) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_10_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_10_n26), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n69), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_10_n27) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_10_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n59), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_10_n25), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_10_n26) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_10_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n69), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_10_n24), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n59), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_10_n30) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_10_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_10_n25), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_10_n24) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_10_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n59), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_10_n25) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_11_U9 ( .A(
        KeyMux_D0_input[11]), .B(KeyMux_D1_input[11]), .S(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_11_n30), .Z(Red_SelectedKey[11]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_11_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_11_n29), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_11_n28), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_11_n27), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_11_n30) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_11_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n75), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_11_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n83), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_11_n27) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_11_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n75), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_11_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n83), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_11_n28) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_11_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_11_n25), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n69), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_11_n26) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_11_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n58), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_11_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_11_n25) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_11_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n69), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_11_n23), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n58), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_11_n29) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_11_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_11_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_11_n23) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_11_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n58), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_11_n24) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_12_U9 ( .A(
        KeyMux_D0_input[12]), .B(KeyMux_D1_input[12]), .S(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_12_n30), .Z(Red_SelectedKey[12]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_12_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_12_n29), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_12_n28), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_12_n27), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_12_n30) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_12_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n75), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_12_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n83), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_12_n27) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_12_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n75), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_12_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n83), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_12_n28) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_12_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_12_n25), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n69), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_12_n26) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_12_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n58), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_12_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_12_n25) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_12_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n69), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_12_n23), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n58), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_12_n29) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_12_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_12_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_12_n23) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_12_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n58), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_12_n24) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_13_U9 ( .A(
        KeyMux_D0_input[13]), .B(KeyMux_D1_input[13]), .S(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_13_n31), .Z(Red_SelectedKey[13]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_13_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_13_n30), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_13_n29), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_13_n28), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_13_n31) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_13_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n75), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_13_n27), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n83), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_13_n28) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_13_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n75), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_13_n27), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n83), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_13_n29) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_13_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_13_n26), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n69), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_13_n27) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_13_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n59), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_13_n25), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_13_n26) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_13_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n69), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_13_n24), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n59), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_13_n30) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_13_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_13_n25), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_13_n24) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_13_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n59), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_13_n25) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_14_U9 ( .A(
        KeyMux_D0_input[14]), .B(KeyMux_D1_input[14]), .S(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_14_n31), .Z(Red_SelectedKey[14]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_14_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_14_n30), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_14_n29), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_14_n28), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_14_n31) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_14_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n75), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_14_n27), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n84), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_14_n28) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_14_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n75), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_14_n27), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n84), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_14_n29) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_14_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_14_n26), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n69), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_14_n27) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_14_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n59), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_14_n25), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_14_n26) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_14_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n69), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_14_n24), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n59), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_14_n30) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_14_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_14_n25), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_14_n24) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_14_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n59), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_14_n25) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_15_U9 ( .A(
        KeyMux_D0_input[15]), .B(KeyMux_D1_input[15]), .S(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_15_n30), .Z(Red_SelectedKey[15]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_15_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_15_n29), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_15_n28), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_15_n27), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_15_n30) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_15_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n74), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_15_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n84), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_15_n27) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_15_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n74), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_15_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n84), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_15_n28) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_15_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_15_n25), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n69), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_15_n26) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_15_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n58), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_15_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_15_n25) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_15_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n69), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_15_n23), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n58), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_15_n29) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_15_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_15_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_15_n23) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_15_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n58), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_15_n24) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_16_U9 ( .A(
        KeyMux_D0_input[16]), .B(KeyMux_D1_input[16]), .S(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_16_n30), .Z(Red_SelectedKey[16]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_16_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_16_n29), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_16_n28), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_16_n27), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_16_n30) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_16_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n78), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_16_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n84), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_16_n27) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_16_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n78), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_16_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n84), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_16_n28) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_16_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_16_n25), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n69), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_16_n26) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_16_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n58), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_16_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_16_n25) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_16_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n69), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_16_n23), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n58), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_16_n29) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_16_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_16_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_16_n23) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_16_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n58), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_16_n24) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_17_U9 ( .A(
        KeyMux_D0_input[17]), .B(KeyMux_D1_input[17]), .S(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_17_n31), .Z(Red_SelectedKey[17]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_17_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_17_n30), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_17_n29), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_17_n28), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_17_n31) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_17_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n76), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_17_n27), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n84), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_17_n28) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_17_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n76), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_17_n27), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n84), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_17_n29) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_17_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_17_n26), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n69), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_17_n27) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_17_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n59), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_17_n25), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_17_n26) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_17_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n69), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_17_n24), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n59), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_17_n30) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_17_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_17_n25), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_17_n24) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_17_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n59), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_17_n25) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_18_U9 ( .A(
        KeyMux_D0_input[18]), .B(KeyMux_D1_input[18]), .S(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_18_n31), .Z(Red_SelectedKey[18]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_18_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_18_n30), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_18_n29), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_18_n28), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_18_n31) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_18_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n75), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_18_n27), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n84), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_18_n28) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_18_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n75), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_18_n27), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n84), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_18_n29) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_18_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_18_n26), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n69), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_18_n27) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_18_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n59), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_18_n25), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_18_n26) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_18_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n69), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_18_n24), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n59), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_18_n30) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_18_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_18_n25), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_18_n24) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_18_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n59), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_18_n25) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_19_U9 ( .A(
        KeyMux_D0_input[19]), .B(KeyMux_D1_input[19]), .S(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_19_n30), .Z(Red_SelectedKey[19]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_19_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_19_n29), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_19_n28), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_19_n27), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_19_n30) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_19_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n76), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_19_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n84), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_19_n27) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_19_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n76), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_19_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n84), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_19_n28) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_19_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_19_n25), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n69), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_19_n26) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_19_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n58), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_19_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_19_n25) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_19_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n69), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_19_n23), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n58), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_19_n29) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_19_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_19_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_19_n23) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_19_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n58), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_19_n24) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_20_U9 ( .A(
        KeyMux_D0_input[20]), .B(KeyMux_D1_input[20]), .S(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_20_n30), .Z(Red_SelectedKey[20]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_20_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_20_n29), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_20_n28), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_20_n27), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_20_n30) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_20_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n75), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_20_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n84), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_20_n27) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_20_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n75), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_20_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n84), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_20_n28) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_20_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_20_n25), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n69), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_20_n26) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_20_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n58), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_20_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_20_n25) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_20_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n69), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_20_n23), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n58), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_20_n29) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_20_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_20_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_20_n23) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_20_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n58), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_20_n24) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_21_U9 ( .A(
        KeyMux_D0_input[21]), .B(KeyMux_D1_input[21]), .S(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_21_n31), .Z(Red_SelectedKey[21]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_21_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_21_n30), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_21_n29), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_21_n28), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_21_n31) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_21_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n76), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_21_n27), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n84), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_21_n28) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_21_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n76), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_21_n27), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n84), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_21_n29) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_21_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_21_n26), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n69), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_21_n27) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_21_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n59), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_21_n25), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_21_n26) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_21_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n69), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_21_n24), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n59), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_21_n30) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_21_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_21_n25), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_21_n24) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_21_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n59), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_21_n25) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_22_U9 ( .A(
        KeyMux_D0_input[22]), .B(KeyMux_D1_input[22]), .S(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_22_n31), .Z(Red_SelectedKey[22]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_22_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_22_n30), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_22_n29), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_22_n28), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_22_n31) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_22_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n76), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_22_n27), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n84), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_22_n28) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_22_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n76), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_22_n27), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n84), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_22_n29) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_22_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_22_n26), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n69), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_22_n27) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_22_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n59), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_22_n25), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_22_n26) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_22_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n69), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_22_n24), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n59), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_22_n30) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_22_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_22_n25), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_22_n24) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_22_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n59), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_22_n25) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_23_U9 ( .A(
        KeyMux_D0_input[23]), .B(KeyMux_D1_input[23]), .S(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_23_n30), .Z(Red_SelectedKey[23]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_23_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_23_n29), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_23_n28), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_23_n27), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_23_n30) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_23_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n76), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_23_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n84), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_23_n27) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_23_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n76), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_23_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n84), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_23_n28) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_23_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_23_n25), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n69), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_23_n26) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_23_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n58), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_23_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_23_n25) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_23_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n69), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_23_n23), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n58), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_23_n29) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_23_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_23_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_23_n23) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_23_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n58), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_23_n24) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_24_U9 ( .A(
        KeyMux_D0_input[24]), .B(KeyMux_D1_input[24]), .S(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_24_n31), .Z(Red_SelectedKey[24]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_24_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_24_n30), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_24_n29), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_24_n28), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_24_n31) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_24_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n76), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_24_n27), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n84), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_24_n28) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_24_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n76), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_24_n27), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n84), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_24_n29) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_24_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_24_n26), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n65), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_24_n27) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_24_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n59), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_24_n25), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_24_n26) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_24_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n65), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_24_n24), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n59), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_24_n30) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_24_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_24_n25), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_24_n24) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_24_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n59), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_24_n25) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_25_U9 ( .A(
        KeyMux_D0_input[25]), .B(KeyMux_D1_input[25]), .S(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_25_n30), .Z(Red_SelectedKey[25]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_25_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_25_n29), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_25_n28), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_25_n27), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_25_n30) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_25_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n76), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_25_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n84), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_25_n27) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_25_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n76), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_25_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n84), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_25_n28) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_25_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_25_n25), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n69), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_25_n26) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_25_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n58), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_25_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_25_n25) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_25_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n69), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_25_n23), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n58), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_25_n29) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_25_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_25_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_25_n23) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_25_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n58), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_25_n24) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_26_U9 ( .A(
        KeyMux_D0_input[26]), .B(KeyMux_D1_input[26]), .S(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_26_n30), .Z(Red_SelectedKey[26]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_26_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_26_n29), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_26_n28), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_26_n27), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_26_n30) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_26_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n75), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_26_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n85), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_26_n27) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_26_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n75), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_26_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n85), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_26_n28) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_26_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_26_n25), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n65), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_26_n26) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_26_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n61), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_26_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_26_n25) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_26_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n65), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_26_n23), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n61), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_26_n29) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_26_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_26_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_26_n23) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_26_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n61), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_26_n24) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_27_U9 ( .A(
        KeyMux_D0_input[27]), .B(KeyMux_D1_input[27]), .S(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_27_n30), .Z(Red_SelectedKey[27]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_27_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_27_n29), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_27_n28), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_27_n27), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_27_n30) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_27_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n76), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_27_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n85), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_27_n27) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_27_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n76), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_27_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n85), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_27_n28) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_27_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_27_n25), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n69), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_27_n26) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_27_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_27_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_27_n25) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_27_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n69), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_27_n23), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_27_n29) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_27_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_27_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_27_n23) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_27_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_27_n24) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_28_U9 ( .A(
        KeyMux_D0_input[28]), .B(KeyMux_D1_input[28]), .S(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_28_n30), .Z(Red_SelectedKey[28]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_28_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_28_n29), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_28_n28), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_28_n27), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_28_n30) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_28_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n75), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_28_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n85), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_28_n27) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_28_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n75), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_28_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n85), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_28_n28) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_28_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_28_n25), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n65), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_28_n26) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_28_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n63), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_28_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_28_n25) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_28_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n65), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_28_n23), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n63), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_28_n29) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_28_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_28_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_28_n23) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_28_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n63), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_28_n24) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_29_U9 ( .A(
        KeyMux_D0_input[29]), .B(KeyMux_D1_input[29]), .S(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_29_n30), .Z(Red_SelectedKey[29]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_29_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_29_n29), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_29_n28), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_29_n27), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_29_n30) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_29_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n76), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_29_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n85), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_29_n27) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_29_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n76), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_29_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n85), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_29_n28) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_29_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_29_n25), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n65), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_29_n26) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_29_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n60), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_29_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_29_n25) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_29_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n65), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_29_n23), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n60), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_29_n29) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_29_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_29_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_29_n23) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_29_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n60), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_29_n24) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_30_U9 ( .A(
        KeyMux_D0_input[30]), .B(KeyMux_D1_input[30]), .S(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_30_n30), .Z(Red_SelectedKey[30]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_30_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_30_n29), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_30_n28), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_30_n27), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_30_n30) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_30_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n76), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_30_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n85), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_30_n27) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_30_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n76), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_30_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n85), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_30_n28) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_30_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_30_n25), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n65), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_30_n26) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_30_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n60), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_30_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_30_n25) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_30_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n65), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_30_n23), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n60), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_30_n29) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_30_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_30_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_30_n23) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_30_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n60), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_30_n24) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_31_U9 ( .A(
        KeyMux_D0_input[31]), .B(KeyMux_D1_input[31]), .S(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_31_n30), .Z(Red_SelectedKey[31]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_31_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_31_n29), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_31_n28), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_31_n27), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_31_n30) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_31_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n76), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_31_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n85), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_31_n27) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_31_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n76), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_31_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n85), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_31_n28) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_31_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_31_n25), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n65), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_31_n26) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_31_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n61), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_31_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_31_n25) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_31_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n65), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_31_n23), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n61), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_31_n29) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_31_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_31_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_31_n23) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_31_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n61), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_31_n24) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_32_U9 ( .A(
        KeyMux_D0_input[32]), .B(KeyMux_D1_input[32]), .S(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_32_n30), .Z(Red_SelectedKey[32]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_32_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_32_n29), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_32_n28), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_32_n27), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_32_n30) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_32_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n76), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_32_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n85), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_32_n27) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_32_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n76), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_32_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n85), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_32_n28) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_32_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_32_n25), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n65), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_32_n26) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_32_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n63), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_32_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_32_n25) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_32_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n65), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_32_n23), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n63), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_32_n29) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_32_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_32_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_32_n23) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_32_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n63), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_32_n24) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_33_U9 ( .A(
        KeyMux_D0_input[33]), .B(KeyMux_D1_input[33]), .S(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_33_n30), .Z(Red_SelectedKey[33]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_33_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_33_n29), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_33_n28), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_33_n27), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_33_n30) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_33_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n76), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_33_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n85), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_33_n27) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_33_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n76), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_33_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n85), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_33_n28) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_33_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_33_n25), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n65), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_33_n26) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_33_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n60), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_33_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_33_n25) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_33_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n65), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_33_n23), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n60), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_33_n29) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_33_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_33_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_33_n23) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_33_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n60), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_33_n24) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_34_U9 ( .A(
        KeyMux_D0_input[34]), .B(KeyMux_D1_input[34]), .S(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_34_n30), .Z(Red_SelectedKey[34]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_34_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_34_n29), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_34_n28), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_34_n27), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_34_n30) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_34_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n76), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_34_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n85), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_34_n27) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_34_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n76), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_34_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n85), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_34_n28) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_34_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_34_n25), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n69), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_34_n26) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_34_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_34_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_34_n25) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_34_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n69), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_34_n23), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_34_n29) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_34_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_34_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_34_n23) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_34_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_34_n24) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_35_U9 ( .A(
        KeyMux_D0_input[35]), .B(KeyMux_D1_input[35]), .S(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_35_n30), .Z(Red_SelectedKey[35]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_35_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_35_n29), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_35_n28), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_35_n27), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_35_n30) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_35_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n76), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_35_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n85), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_35_n27) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_35_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n76), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_35_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n85), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_35_n28) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_35_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_35_n25), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n69), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_35_n26) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_35_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n63), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_35_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_35_n25) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_35_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n69), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_35_n23), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n63), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_35_n29) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_35_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_35_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_35_n23) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_35_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n63), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_35_n24) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_36_U9 ( .A(
        KeyMux_D0_input[36]), .B(KeyMux_D1_input[36]), .S(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_36_n30), .Z(Red_SelectedKey[36]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_36_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_36_n29), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_36_n28), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_36_n27), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_36_n30) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_36_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n76), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_36_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n85), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_36_n27) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_36_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n76), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_36_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n85), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_36_n28) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_36_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_36_n25), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n69), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_36_n26) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_36_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n60), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_36_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_36_n25) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_36_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n69), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_36_n23), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n60), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_36_n29) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_36_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_36_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_36_n23) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_36_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n60), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_36_n24) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_37_U9 ( .A(
        KeyMux_D0_input[37]), .B(KeyMux_D1_input[37]), .S(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_37_n30), .Z(Red_SelectedKey[37]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_37_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_37_n29), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_37_n28), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_37_n27), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_37_n30) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_37_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n76), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_37_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n85), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_37_n27) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_37_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n76), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_37_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n85), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_37_n28) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_37_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_37_n25), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n69), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_37_n26) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_37_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_37_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_37_n25) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_37_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n69), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_37_n23), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_37_n29) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_37_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_37_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_37_n23) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_37_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_37_n24) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_38_U9 ( .A(
        KeyMux_D0_input[38]), .B(KeyMux_D1_input[38]), .S(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_38_n30), .Z(Red_SelectedKey[38]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_38_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_38_n29), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_38_n28), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_38_n27), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_38_n30) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_38_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n77), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_38_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n86), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_38_n27) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_38_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n77), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_38_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n86), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_38_n28) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_38_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_38_n25), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n70), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_38_n26) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_38_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_38_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_38_n25) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_38_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n70), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_38_n23), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_38_n29) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_38_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_38_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_38_n23) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_38_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_38_n24) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_39_U9 ( .A(
        KeyMux_D0_input[39]), .B(KeyMux_D1_input[39]), .S(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_39_n30), .Z(Red_SelectedKey[39]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_39_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_39_n29), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_39_n28), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_39_n27), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_39_n30) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_39_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n77), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_39_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n86), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_39_n27) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_39_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n77), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_39_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n86), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_39_n28) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_39_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_39_n25), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n70), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_39_n26) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_39_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_39_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_39_n25) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_39_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n70), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_39_n23), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_39_n29) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_39_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_39_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_39_n23) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_39_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_39_n24) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_40_U9 ( .A(
        KeyMux_D0_input[40]), .B(KeyMux_D1_input[40]), .S(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_40_n30), .Z(Red_SelectedKey[40]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_40_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_40_n29), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_40_n28), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_40_n27), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_40_n30) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_40_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n77), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_40_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n86), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_40_n27) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_40_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n77), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_40_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n86), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_40_n28) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_40_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_40_n25), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n70), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_40_n26) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_40_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_40_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_40_n25) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_40_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n70), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_40_n23), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_40_n29) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_40_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_40_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_40_n23) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_40_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_40_n24) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_41_U9 ( .A(
        KeyMux_D0_input[41]), .B(KeyMux_D1_input[41]), .S(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_41_n30), .Z(Red_SelectedKey[41]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_41_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_41_n29), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_41_n28), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_41_n27), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_41_n30) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_41_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n77), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_41_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n86), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_41_n27) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_41_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n77), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_41_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n86), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_41_n28) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_41_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_41_n25), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n70), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_41_n26) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_41_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_41_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_41_n25) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_41_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n70), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_41_n23), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_41_n29) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_41_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_41_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_41_n23) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_41_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_41_n24) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_42_U9 ( .A(
        KeyMux_D0_input[42]), .B(KeyMux_D1_input[42]), .S(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_42_n30), .Z(Red_SelectedKey[42]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_42_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_42_n29), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_42_n28), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_42_n27), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_42_n30) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_42_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n77), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_42_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n86), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_42_n27) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_42_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n77), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_42_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n86), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_42_n28) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_42_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_42_n25), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n70), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_42_n26) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_42_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_42_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_42_n25) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_42_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n70), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_42_n23), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_42_n29) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_42_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_42_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_42_n23) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_42_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_42_n24) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_43_U9 ( .A(
        KeyMux_D0_input[43]), .B(KeyMux_D1_input[43]), .S(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_43_n30), .Z(Red_SelectedKey[43]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_43_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_43_n29), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_43_n28), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_43_n27), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_43_n30) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_43_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n77), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_43_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n86), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_43_n27) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_43_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n77), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_43_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n86), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_43_n28) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_43_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_43_n25), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n70), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_43_n26) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_43_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_43_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_43_n25) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_43_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n70), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_43_n23), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_43_n29) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_43_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_43_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_43_n23) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_43_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_43_n24) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_44_U9 ( .A(
        KeyMux_D0_input[44]), .B(KeyMux_D1_input[44]), .S(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_44_n30), .Z(Red_SelectedKey[44]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_44_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_44_n29), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_44_n28), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_44_n27), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_44_n30) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_44_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n77), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_44_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n86), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_44_n27) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_44_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n77), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_44_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n86), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_44_n28) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_44_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_44_n25), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n70), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_44_n26) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_44_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_44_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_44_n25) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_44_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n70), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_44_n23), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_44_n29) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_44_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_44_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_44_n23) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_44_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_44_n24) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_45_U9 ( .A(
        KeyMux_D0_input[45]), .B(KeyMux_D1_input[45]), .S(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_45_n30), .Z(Red_SelectedKey[45]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_45_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_45_n29), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_45_n28), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_45_n27), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_45_n30) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_45_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n77), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_45_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n86), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_45_n27) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_45_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n77), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_45_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n86), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_45_n28) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_45_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_45_n25), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n70), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_45_n26) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_45_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_45_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_45_n25) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_45_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n70), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_45_n23), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_45_n29) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_45_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_45_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_45_n23) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_45_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_45_n24) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_46_U9 ( .A(
        KeyMux_D0_input[46]), .B(KeyMux_D1_input[46]), .S(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_46_n31), .Z(Red_SelectedKey[46]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_46_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_46_n30), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_46_n29), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_46_n28), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_46_n31) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_46_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n77), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_46_n27), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n86), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_46_n28) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_46_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n77), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_46_n27), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n86), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_46_n29) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_46_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_46_n26), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n70), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_46_n27) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_46_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n59), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_46_n25), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_46_n26) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_46_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n70), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_46_n24), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n59), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_46_n30) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_46_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_46_n25), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_46_n24) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_46_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n59), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_46_n25) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_47_U9 ( .A(
        KeyMux_D0_input[47]), .B(KeyMux_D1_input[47]), .S(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_47_n30), .Z(Red_SelectedKey[47]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_47_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_47_n29), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_47_n28), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_47_n27), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_47_n30) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_47_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n77), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_47_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n86), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_47_n27) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_47_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n77), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_47_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n86), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_47_n28) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_47_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_47_n25), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n70), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_47_n26) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_47_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_47_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_47_n25) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_47_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n70), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_47_n23), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_47_n29) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_47_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_47_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_47_n23) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_47_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_47_n24) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_48_U9 ( .A(
        KeyMux_D0_input[48]), .B(KeyMux_D1_input[48]), .S(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_48_n30), .Z(Red_SelectedKey[48]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_48_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_48_n29), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_48_n28), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_48_n27), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_48_n30) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_48_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n77), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_48_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n86), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_48_n27) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_48_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n77), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_48_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n86), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_48_n28) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_48_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_48_n25), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n70), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_48_n26) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_48_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_48_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_48_n25) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_48_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n70), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_48_n23), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_48_n29) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_48_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_48_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_48_n23) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_48_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_48_n24) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_49_U9 ( .A(
        KeyMux_D0_input[49]), .B(KeyMux_D1_input[49]), .S(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_49_n30), .Z(Red_SelectedKey[49]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_49_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_49_n29), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_49_n28), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_49_n27), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_49_n30) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_49_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n77), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_49_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n86), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_49_n27) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_49_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n77), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_49_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n86), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_49_n28) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_49_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_49_n25), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n70), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_49_n26) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_49_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_49_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_49_n25) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_49_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n70), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_49_n23), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_49_n29) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_49_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_49_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_49_n23) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_49_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_49_n24) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_50_U9 ( .A(
        KeyMux_D0_input[50]), .B(KeyMux_D1_input[50]), .S(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_50_n30), .Z(Red_SelectedKey[50]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_50_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_50_n29), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_50_n28), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_50_n27), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_50_n30) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_50_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n77), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_50_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n89), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_50_n27) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_50_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n77), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_50_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n89), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_50_n28) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_50_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_50_n25), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n66), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_50_n26) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_50_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n60), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_50_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_50_n25) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_50_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n66), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_50_n23), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n60), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_50_n29) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_50_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_50_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_50_n23) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_50_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n60), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_50_n24) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_51_U9 ( .A(
        KeyMux_D0_input[51]), .B(KeyMux_D1_input[51]), .S(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_51_n30), .Z(Red_SelectedKey[51]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_51_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_51_n29), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_51_n28), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_51_n27), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_51_n30) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_51_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n78), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_51_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n84), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_51_n27) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_51_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n78), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_51_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n84), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_51_n28) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_51_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_51_n25), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n66), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_51_n26) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_51_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n63), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_51_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_51_n25) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_51_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n66), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_51_n23), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n63), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_51_n29) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_51_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_51_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_51_n23) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_51_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n63), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_51_n24) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_52_U9 ( .A(
        KeyMux_D0_input[52]), .B(KeyMux_D1_input[52]), .S(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_52_n30), .Z(Red_SelectedKey[52]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_52_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_52_n29), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_52_n28), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_52_n27), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_52_n30) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_52_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n78), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_52_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n89), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_52_n27) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_52_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n78), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_52_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n89), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_52_n28) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_52_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_52_n25), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n66), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_52_n26) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_52_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n63), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_52_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_52_n25) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_52_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n66), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_52_n23), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n63), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_52_n29) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_52_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_52_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_52_n23) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_52_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n63), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_52_n24) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_53_U9 ( .A(
        KeyMux_D0_input[53]), .B(KeyMux_D1_input[53]), .S(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_53_n30), .Z(Red_SelectedKey[53]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_53_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_53_n29), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_53_n28), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_53_n27), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_53_n30) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_53_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n78), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_53_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n84), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_53_n27) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_53_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n78), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_53_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n84), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_53_n28) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_53_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_53_n25), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n66), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_53_n26) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_53_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n60), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_53_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_53_n25) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_53_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n66), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_53_n23), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n60), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_53_n29) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_53_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_53_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_53_n23) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_53_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n60), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_53_n24) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_54_U9 ( .A(
        KeyMux_D0_input[54]), .B(KeyMux_D1_input[54]), .S(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_54_n30), .Z(Red_SelectedKey[54]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_54_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_54_n29), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_54_n28), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_54_n27), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_54_n30) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_54_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n78), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_54_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n84), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_54_n27) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_54_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n78), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_54_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n84), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_54_n28) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_54_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_54_n25), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n70), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_54_n26) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_54_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n60), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_54_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_54_n25) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_54_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n70), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_54_n23), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n60), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_54_n29) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_54_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_54_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_54_n23) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_54_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n60), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_54_n24) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_55_U9 ( .A(
        KeyMux_D0_input[55]), .B(KeyMux_D1_input[55]), .S(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_55_n30), .Z(Red_SelectedKey[55]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_55_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_55_n29), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_55_n28), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_55_n27), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_55_n30) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_55_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n78), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_55_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n89), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_55_n27) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_55_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n78), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_55_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n89), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_55_n28) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_55_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_55_n25), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n70), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_55_n26) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_55_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n63), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_55_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_55_n25) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_55_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n70), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_55_n23), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n63), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_55_n29) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_55_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_55_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_55_n23) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_55_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n63), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_55_n24) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_56_U9 ( .A(
        KeyMux_D0_input[56]), .B(KeyMux_D1_input[56]), .S(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_56_n30), .Z(Red_SelectedKey[56]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_56_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_56_n29), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_56_n28), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_56_n27), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_56_n30) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_56_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n80), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_56_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n87), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_56_n27) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_56_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n80), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_56_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n87), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_56_n28) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_56_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_56_n25), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n67), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_56_n26) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_56_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n63), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_56_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_56_n25) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_56_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n67), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_56_n23), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n63), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_56_n29) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_56_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_56_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_56_n23) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_56_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n63), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_56_n24) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_57_U9 ( .A(
        KeyMux_D0_input[57]), .B(KeyMux_D1_input[57]), .S(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_57_n31), .Z(Red_SelectedKey[57]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_57_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_57_n30), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_57_n29), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_57_n28), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_57_n31) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_57_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n80), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_57_n27), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n86), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_57_n28) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_57_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n80), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_57_n27), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n86), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_57_n29) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_57_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_57_n26), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n67), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_57_n27) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_57_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n59), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_57_n25), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_57_n26) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_57_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n67), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_57_n24), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n59), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_57_n30) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_57_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_57_n25), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_57_n24) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_57_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n59), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_57_n25) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_58_U9 ( .A(
        KeyMux_D0_input[58]), .B(KeyMux_D1_input[58]), .S(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_58_n30), .Z(Red_SelectedKey[58]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_58_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_58_n29), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_58_n28), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_58_n27), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_58_n30) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_58_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n80), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_58_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n87), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_58_n27) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_58_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n80), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_58_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n87), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_58_n28) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_58_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_58_n25), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n67), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_58_n26) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_58_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n60), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_58_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_58_n25) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_58_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n67), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_58_n23), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n60), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_58_n29) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_58_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_58_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_58_n23) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_58_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n60), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_58_n24) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_59_U9 ( .A(
        KeyMux_D0_input[59]), .B(KeyMux_D1_input[59]), .S(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_59_n30), .Z(Red_SelectedKey[59]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_59_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_59_n29), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_59_n28), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_59_n27), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_59_n30) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_59_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n80), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_59_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n86), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_59_n27) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_59_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n80), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_59_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n86), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_59_n28) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_59_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_59_n25), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n67), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_59_n26) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_59_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n63), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_59_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_59_n25) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_59_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n67), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_59_n23), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n63), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_59_n29) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_59_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_59_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_59_n23) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_59_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n63), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_59_n24) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_60_U9 ( .A(
        KeyMux_D0_input[60]), .B(KeyMux_D1_input[60]), .S(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_60_n30), .Z(Red_SelectedKey[60]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_60_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_60_n29), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_60_n28), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_60_n27), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_60_n30) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_60_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n80), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_60_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n87), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_60_n27) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_60_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n80), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_60_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n87), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_60_n28) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_60_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_60_n25), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n67), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_60_n26) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_60_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n58), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_60_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_60_n25) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_60_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n67), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_60_n23), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n58), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_60_n29) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_60_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_60_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_60_n23) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_60_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n58), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_60_n24) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_61_U9 ( .A(
        KeyMux_D0_input[61]), .B(KeyMux_D1_input[61]), .S(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_61_n30), .Z(Red_SelectedKey[61]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_61_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_61_n29), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_61_n28), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_61_n27), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_61_n30) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_61_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n80), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_61_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n86), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_61_n27) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_61_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n80), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_61_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n86), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_61_n28) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_61_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_61_n25), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n67), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_61_n26) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_61_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n63), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_61_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_61_n25) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_61_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n67), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_61_n23), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n63), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_61_n29) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_61_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_61_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_61_n23) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_61_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n63), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_61_n24) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_62_U9 ( .A(
        KeyMux_D0_input[62]), .B(KeyMux_D1_input[62]), .S(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_62_n30), .Z(Red_SelectedKey[62]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_62_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_62_n29), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_62_n28), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_62_n27), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_62_n30) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_62_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n80), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_62_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n87), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_62_n27) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_62_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n80), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_62_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n87), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_62_n28) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_62_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_62_n25), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n67), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_62_n26) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_62_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_62_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_62_n25) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_62_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n67), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_62_n23), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_62_n29) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_62_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_62_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_62_n23) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_62_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_62_n24) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_63_U9 ( .A(
        KeyMux_D0_input[63]), .B(KeyMux_D1_input[63]), .S(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_63_n31), .Z(Red_SelectedKey[63]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_63_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_63_n30), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_63_n29), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_63_n28), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_63_n31) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_63_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n80), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_63_n27), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n86), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_63_n28) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_63_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n80), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_63_n27), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n86), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_63_n29) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_63_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_63_n26), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n67), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_63_n27) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_63_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n59), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_63_n25), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_63_n26) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_63_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n67), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_63_n24), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n59), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_63_n30) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_63_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_63_n25), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_63_n24) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_63_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n59), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_63_n25) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_64_U9 ( .A(
        KeyMux_D0_input[64]), .B(KeyMux_D1_input[64]), .S(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_64_n30), .Z(Red_SelectedKey[64]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_64_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_64_n29), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_64_n28), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_64_n27), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_64_n30) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_64_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n80), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_64_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n87), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_64_n27) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_64_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n80), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_64_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n87), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_64_n28) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_64_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_64_n25), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n71), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_64_n26) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_64_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_64_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_64_n25) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_64_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n71), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_64_n23), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_64_n29) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_64_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_64_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_64_n23) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_64_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_64_n24) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_65_U9 ( .A(
        KeyMux_D0_input[65]), .B(KeyMux_D1_input[65]), .S(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_65_n30), .Z(Red_SelectedKey[65]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_65_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_65_n29), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_65_n28), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_65_n27), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_65_n30) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_65_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n80), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_65_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n86), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_65_n27) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_65_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n80), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_65_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n86), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_65_n28) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_65_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_65_n25), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n71), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_65_n26) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_65_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n61), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_65_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_65_n25) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_65_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n71), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_65_n23), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n61), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_65_n29) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_65_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_65_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_65_n23) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_65_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n61), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_65_n24) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_66_U9 ( .A(
        KeyMux_D0_input[66]), .B(KeyMux_D1_input[66]), .S(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_66_n30), .Z(Red_SelectedKey[66]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_66_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_66_n29), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_66_n28), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_66_n27), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_66_n30) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_66_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n80), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_66_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n87), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_66_n27) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_66_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n80), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_66_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n87), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_66_n28) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_66_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_66_n25), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n71), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_66_n26) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_66_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_66_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_66_n25) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_66_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n71), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_66_n23), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_66_n29) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_66_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_66_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_66_n23) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_66_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_66_n24) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_67_U9 ( .A(
        KeyMux_D0_input[67]), .B(KeyMux_D1_input[67]), .S(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_67_n30), .Z(Red_SelectedKey[67]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_67_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_67_n29), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_67_n28), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_67_n27), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_67_n30) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_67_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n80), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_67_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n86), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_67_n27) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_67_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n80), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_67_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n86), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_67_n28) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_67_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_67_n25), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n71), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_67_n26) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_67_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_67_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_67_n25) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_67_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n71), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_67_n23), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_67_n29) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_67_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_67_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_67_n23) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_67_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_67_n24) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_68_U9 ( .A(
        KeyMux_D0_input[68]), .B(KeyMux_D1_input[68]), .S(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_68_n30), .Z(Red_SelectedKey[68]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_68_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_68_n29), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_68_n28), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_68_n27), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_68_n30) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_68_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n80), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_68_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n87), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_68_n27) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_68_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n80), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_68_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n87), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_68_n28) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_68_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_68_n25), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n71), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_68_n26) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_68_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_68_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_68_n25) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_68_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n71), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_68_n23), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_68_n29) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_68_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_68_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_68_n23) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_68_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_68_n24) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_69_U9 ( .A(
        KeyMux_D0_input[69]), .B(KeyMux_D1_input[69]), .S(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_69_n30), .Z(Red_SelectedKey[69]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_69_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_69_n29), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_69_n28), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_69_n27), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_69_n30) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_69_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n80), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_69_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n86), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_69_n27) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_69_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n80), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_69_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n86), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_69_n28) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_69_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_69_n25), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n71), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_69_n26) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_69_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_69_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_69_n25) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_69_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n71), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_69_n23), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_69_n29) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_69_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_69_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_69_n23) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_69_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_69_n24) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_70_U9 ( .A(
        KeyMux_D0_input[70]), .B(KeyMux_D1_input[70]), .S(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_70_n30), .Z(Red_SelectedKey[70]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_70_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_70_n29), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_70_n28), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_70_n27), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_70_n30) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_70_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n79), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_70_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n84), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_70_n27) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_70_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n79), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_70_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n84), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_70_n28) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_70_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_70_n25), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n71), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_70_n26) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_70_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_70_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_70_n25) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_70_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n71), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_70_n23), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_70_n29) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_70_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_70_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_70_n23) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_70_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_70_n24) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_71_U9 ( .A(
        KeyMux_D0_input[71]), .B(KeyMux_D1_input[71]), .S(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_71_n30), .Z(Red_SelectedKey[71]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_71_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_71_n29), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_71_n28), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_71_n27), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_71_n30) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_71_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n74), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_71_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n89), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_71_n27) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_71_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n74), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_71_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n89), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_71_n28) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_71_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_71_n25), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n71), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_71_n26) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_71_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_71_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_71_n25) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_71_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n71), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_71_n23), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_71_n29) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_71_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_71_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_71_n23) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_71_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_71_n24) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_72_U9 ( .A(
        KeyMux_D0_input[72]), .B(KeyMux_D1_input[72]), .S(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_72_n30), .Z(Red_SelectedKey[72]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_72_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_72_n29), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_72_n28), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_72_n27), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_72_n30) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_72_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n79), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_72_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n85), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_72_n27) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_72_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n79), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_72_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n85), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_72_n28) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_72_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_72_n25), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n71), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_72_n26) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_72_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_72_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_72_n25) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_72_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n71), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_72_n23), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_72_n29) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_72_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_72_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_72_n23) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_72_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_72_n24) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_73_U9 ( .A(
        KeyMux_D0_input[73]), .B(KeyMux_D1_input[73]), .S(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_73_n30), .Z(Red_SelectedKey[73]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_73_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_73_n29), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_73_n28), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_73_n27), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_73_n30) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_73_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n80), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_73_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n83), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_73_n27) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_73_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n80), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_73_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n83), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_73_n28) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_73_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_73_n25), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n71), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_73_n26) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_73_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_73_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_73_n25) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_73_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n71), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_73_n23), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_73_n29) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_73_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_73_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_73_n23) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_73_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_73_n24) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_74_U9 ( .A(
        KeyMux_D0_input[74]), .B(KeyMux_D1_input[74]), .S(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_74_n30), .Z(Red_SelectedKey[74]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_74_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_74_n29), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_74_n28), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_74_n27), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_74_n30) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_74_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n79), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_74_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n85), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_74_n27) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_74_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n79), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_74_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n85), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_74_n28) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_74_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_74_n25), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n71), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_74_n26) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_74_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_74_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_74_n25) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_74_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n71), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_74_n23), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_74_n29) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_74_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_74_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_74_n23) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_74_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_74_n24) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_75_U9 ( .A(
        KeyMux_D0_input[75]), .B(KeyMux_D1_input[75]), .S(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_75_n30), .Z(Red_SelectedKey[75]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_75_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_75_n29), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_75_n28), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_75_n27), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_75_n30) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_75_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n79), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_75_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n88), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_75_n27) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_75_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n79), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_75_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n88), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_75_n28) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_75_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_75_n25), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n71), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_75_n26) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_75_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_75_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_75_n25) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_75_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n71), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_75_n23), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_75_n29) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_75_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_75_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_75_n23) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_75_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_75_n24) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_76_U9 ( .A(
        KeyMux_D0_input[76]), .B(KeyMux_D1_input[76]), .S(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_76_n30), .Z(Red_SelectedKey[76]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_76_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_76_n29), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_76_n28), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_76_n27), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_76_n30) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_76_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n79), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_76_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n89), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_76_n27) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_76_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n79), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_76_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n89), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_76_n28) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_76_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_76_n25), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n71), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_76_n26) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_76_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_76_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_76_n25) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_76_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n71), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_76_n23), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_76_n29) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_76_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_76_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_76_n23) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_76_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_76_n24) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_77_U9 ( .A(
        KeyMux_D0_input[77]), .B(KeyMux_D1_input[77]), .S(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_77_n30), .Z(Red_SelectedKey[77]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_77_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_77_n29), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_77_n28), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_77_n27), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_77_n30) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_77_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n79), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_77_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n88), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_77_n27) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_77_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n79), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_77_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n88), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_77_n28) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_77_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_77_n25), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n71), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_77_n26) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_77_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_77_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_77_n25) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_77_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n71), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_77_n23), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_77_n29) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_77_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_77_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_77_n23) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_77_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_77_n24) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_78_U9 ( .A(
        KeyMux_D0_input[78]), .B(KeyMux_D1_input[78]), .S(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_78_n30), .Z(Red_SelectedKey[78]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_78_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_78_n29), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_78_n28), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_78_n27), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_78_n30) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_78_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n81), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_78_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n88), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_78_n27) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_78_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n81), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_78_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n88), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_78_n28) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_78_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_78_n25), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n69), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_78_n26) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_78_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n61), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_78_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_78_n25) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_78_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n69), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_78_n23), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n61), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_78_n29) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_78_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_78_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_78_n23) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_78_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n61), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_78_n24) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_79_U9 ( .A(
        KeyMux_D0_input[79]), .B(KeyMux_D1_input[79]), .S(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_79_n30), .Z(Red_SelectedKey[79]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_79_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_79_n29), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_79_n28), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_79_n27), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_79_n30) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_79_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n81), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_79_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n88), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_79_n27) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_79_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n81), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_79_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n88), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_79_n28) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_79_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_79_n25), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n71), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_79_n26) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_79_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n61), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_79_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_79_n25) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_79_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n71), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_79_n23), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n61), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_79_n29) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_79_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_79_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_79_n23) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_79_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n61), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_79_n24) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_80_U9 ( .A(
        KeyMux_D0_input[80]), .B(KeyMux_D1_input[80]), .S(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_80_n30), .Z(Red_SelectedKey[80]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_80_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_80_n29), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_80_n28), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_80_n27), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_80_n30) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_80_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n81), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_80_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n88), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_80_n27) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_80_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n81), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_80_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n88), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_80_n28) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_80_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_80_n25), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n71), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_80_n26) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_80_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n61), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_80_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_80_n25) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_80_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n71), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_80_n23), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n61), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_80_n29) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_80_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_80_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_80_n23) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_80_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n61), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_80_n24) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_81_U9 ( .A(
        KeyMux_D0_input[81]), .B(KeyMux_D1_input[81]), .S(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_81_n30), .Z(Red_SelectedKey[81]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_81_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_81_n29), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_81_n28), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_81_n27), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_81_n30) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_81_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n81), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_81_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n88), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_81_n27) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_81_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n81), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_81_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n88), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_81_n28) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_81_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_81_n25), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n70), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_81_n26) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_81_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n61), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_81_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_81_n25) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_81_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n70), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_81_n23), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n61), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_81_n29) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_81_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_81_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_81_n23) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_81_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n61), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_81_n24) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_82_U9 ( .A(
        KeyMux_D0_input[82]), .B(KeyMux_D1_input[82]), .S(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_82_n30), .Z(Red_SelectedKey[82]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_82_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_82_n29), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_82_n28), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_82_n27), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_82_n30) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_82_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n81), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_82_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n88), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_82_n27) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_82_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n81), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_82_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n88), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_82_n28) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_82_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_82_n25), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n70), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_82_n26) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_82_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n61), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_82_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_82_n25) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_82_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n70), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_82_n23), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n61), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_82_n29) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_82_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_82_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_82_n23) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_82_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n61), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_82_n24) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_83_U9 ( .A(
        KeyMux_D0_input[83]), .B(KeyMux_D1_input[83]), .S(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_83_n30), .Z(Red_SelectedKey[83]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_83_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_83_n29), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_83_n28), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_83_n27), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_83_n30) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_83_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n81), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_83_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n88), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_83_n27) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_83_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n81), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_83_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n88), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_83_n28) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_83_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_83_n25), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n69), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_83_n26) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_83_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n61), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_83_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_83_n25) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_83_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n69), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_83_n23), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n61), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_83_n29) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_83_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_83_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_83_n23) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_83_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n61), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_83_n24) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_84_U9 ( .A(
        KeyMux_D0_input[84]), .B(KeyMux_D1_input[84]), .S(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_84_n30), .Z(Red_SelectedKey[84]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_84_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_84_n29), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_84_n28), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_84_n27), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_84_n30) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_84_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n81), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_84_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n88), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_84_n27) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_84_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n81), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_84_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n88), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_84_n28) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_84_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_84_n25), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n70), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_84_n26) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_84_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n61), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_84_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_84_n25) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_84_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n70), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_84_n23), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n61), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_84_n29) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_84_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_84_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_84_n23) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_84_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n61), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_84_n24) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_85_U9 ( .A(
        KeyMux_D0_input[85]), .B(KeyMux_D1_input[85]), .S(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_85_n30), .Z(Red_SelectedKey[85]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_85_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_85_n29), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_85_n28), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_85_n27), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_85_n30) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_85_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n81), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_85_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n88), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_85_n27) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_85_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n81), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_85_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n88), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_85_n28) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_85_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_85_n25), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n69), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_85_n26) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_85_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n61), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_85_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_85_n25) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_85_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n69), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_85_n23), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n61), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_85_n29) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_85_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_85_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_85_n23) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_85_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n61), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_85_n24) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_86_U9 ( .A(
        KeyMux_D0_input[86]), .B(KeyMux_D1_input[86]), .S(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_86_n30), .Z(Red_SelectedKey[86]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_86_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_86_n29), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_86_n28), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_86_n27), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_86_n30) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_86_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n81), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_86_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n88), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_86_n27) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_86_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n81), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_86_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n88), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_86_n28) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_86_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_86_n25), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n71), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_86_n26) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_86_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n61), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_86_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_86_n25) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_86_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n71), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_86_n23), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n61), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_86_n29) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_86_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_86_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_86_n23) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_86_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n61), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_86_n24) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_87_U9 ( .A(
        KeyMux_D0_input[87]), .B(KeyMux_D1_input[87]), .S(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_87_n31), .Z(Red_SelectedKey[87]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_87_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_87_n30), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_87_n29), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_87_n28), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_87_n31) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_87_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n81), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_87_n27), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n88), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_87_n28) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_87_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n81), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_87_n27), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n88), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_87_n29) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_87_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_87_n26), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n70), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_87_n27) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_87_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n59), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_87_n25), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_87_n26) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_87_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n70), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_87_n24), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n59), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_87_n30) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_87_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_87_n25), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_87_n24) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_87_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n59), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_87_n25) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_88_U9 ( .A(
        KeyMux_D0_input[88]), .B(KeyMux_D1_input[88]), .S(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_88_n31), .Z(Red_SelectedKey[88]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_88_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_88_n30), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_88_n29), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_88_n28), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_88_n31) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_88_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n81), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_88_n27), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n88), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_88_n28) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_88_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n81), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_88_n27), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n88), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_88_n29) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_88_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_88_n26), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n69), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_88_n27) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_88_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n59), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_88_n25), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_88_n26) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_88_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n69), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_88_n24), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n59), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_88_n30) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_88_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_88_n25), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_88_n24) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_88_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n59), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_88_n25) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_89_U9 ( .A(
        KeyMux_D0_input[89]), .B(KeyMux_D1_input[89]), .S(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_89_n31), .Z(Red_SelectedKey[89]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_89_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_89_n30), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_89_n29), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_89_n28), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_89_n31) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_89_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n81), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_89_n27), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n88), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_89_n28) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_89_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n81), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_89_n27), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n88), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_89_n29) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_89_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_89_n26), .B(n3), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_89_n27) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_89_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n59), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_89_n25), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_89_n26) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_89_U3 ( .A1(n3), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_89_n24), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n59), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_89_n30) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_89_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_89_n25), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_89_n24) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_89_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n59), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_89_n25) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_90_U9 ( .A(
        KeyMux_D0_input[90]), .B(KeyMux_D1_input[90]), .S(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_90_n31), .Z(Red_SelectedKey[90]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_90_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_90_n30), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_90_n29), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_90_n28), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_90_n31) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_90_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n81), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_90_n27), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n86), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_90_n28) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_90_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n81), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_90_n27), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n86), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_90_n29) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_90_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_90_n26), .B(n3), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_90_n27) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_90_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_90_n25), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_90_n26) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_90_U3 ( .A1(n3), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_90_n24), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_90_n30) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_90_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_90_n25), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_90_n24) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_90_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_90_n25) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_91_U9 ( .A(
        KeyMux_D0_input[91]), .B(KeyMux_D1_input[91]), .S(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_91_n31), .Z(Red_SelectedKey[91]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_91_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_91_n30), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_91_n29), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_91_n28), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_91_n31) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_91_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n82), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_91_n27), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n87), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_91_n28) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_91_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n82), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_91_n27), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n87), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_91_n29) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_91_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_91_n26), .B(n3), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_91_n27) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_91_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n58), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_91_n25), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_91_n26) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_91_U3 ( .A1(n3), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_91_n24), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n58), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_91_n30) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_91_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_91_n25), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_91_n24) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_91_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n58), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_91_n25) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_92_U9 ( .A(
        KeyMux_D0_input[92]), .B(KeyMux_D1_input[92]), .S(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_92_n31), .Z(Red_SelectedKey[92]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_92_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_92_n30), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_92_n29), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_92_n28), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_92_n31) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_92_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n82), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_92_n27), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n86), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_92_n28) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_92_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n82), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_92_n27), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n86), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_92_n29) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_92_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_92_n26), .B(n3), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_92_n27) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_92_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n58), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_92_n25), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_92_n26) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_92_U3 ( .A1(n3), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_92_n24), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n58), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_92_n30) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_92_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_92_n25), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_92_n24) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_92_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n58), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_92_n25) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_93_U9 ( .A(
        KeyMux_D0_input[93]), .B(KeyMux_D1_input[93]), .S(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_93_n31), .Z(Red_SelectedKey[93]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_93_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_93_n30), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_93_n29), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_93_n28), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_93_n31) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_93_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n81), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_93_n27), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n86), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_93_n28) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_93_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n81), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_93_n27), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n86), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_93_n29) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_93_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_93_n26), .B(n3), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_93_n27) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_93_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_93_n25), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_93_n26) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_93_U3 ( .A1(n3), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_93_n24), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_93_n30) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_93_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_93_n25), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_93_n24) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_93_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_93_n25) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_94_U9 ( .A(
        KeyMux_D0_input[94]), .B(KeyMux_D1_input[94]), .S(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_94_n31), .Z(Red_SelectedKey[94]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_94_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_94_n30), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_94_n29), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_94_n28), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_94_n31) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_94_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n82), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_94_n27), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n87), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_94_n28) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_94_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n82), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_94_n27), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n87), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_94_n29) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_94_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_94_n26), .B(n3), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_94_n27) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_94_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n63), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_94_n25), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_94_n26) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_94_U3 ( .A1(n3), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_94_n24), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n63), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_94_n30) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_94_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_94_n25), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_94_n24) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_94_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n63), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_94_n25) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_95_U9 ( .A(
        KeyMux_D0_input[95]), .B(KeyMux_D1_input[95]), .S(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_95_n32), .Z(Red_SelectedKey[95]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_95_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_95_n31), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_95_n30), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_95_n29), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_95_n32) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_95_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n81), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_95_n28), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n87), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_95_n29) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_95_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n81), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_95_n28), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n87), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_95_n30) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_95_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_95_n27), .B(n3), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_95_n28) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_95_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n59), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_95_n26), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_95_n27) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_95_U3 ( .A1(n3), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_95_n25), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n59), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_95_n31) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_95_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_95_n26), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_95_n25) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_95_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n59), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_95_n26) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_96_U9 ( .A(
        KeyMux_D0_input[96]), .B(KeyMux_D1_input[96]), .S(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_96_n32), .Z(Red_SelectedKey[96]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_96_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_96_n31), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_96_n30), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_96_n29), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_96_n32) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_96_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n82), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_96_n28), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n86), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_96_n29) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_96_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n82), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_96_n28), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n86), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_96_n30) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_96_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_96_n27), .B(n3), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_96_n28) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_96_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n59), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_96_n26), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_96_n27) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_96_U3 ( .A1(n3), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_96_n25), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n59), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_96_n31) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_96_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_96_n26), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_96_n25) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_96_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n59), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_96_n26) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_97_U9 ( .A(
        KeyMux_D0_input[97]), .B(KeyMux_D1_input[97]), .S(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_97_n30), .Z(Red_SelectedKey[97]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_97_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_97_n29), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_97_n28), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_97_n27), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_97_n30) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_97_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n82), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_97_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n87), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_97_n27) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_97_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n82), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_97_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n87), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_97_n28) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_97_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_97_n25), .B(n3), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_97_n26) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_97_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n60), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_97_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_97_n25) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_97_U3 ( .A1(n3), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_97_n23), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n60), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_97_n29) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_97_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_97_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_97_n23) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_97_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n60), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_97_n24) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_98_U9 ( .A(
        KeyMux_D0_input[98]), .B(KeyMux_D1_input[98]), .S(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_98_n30), .Z(Red_SelectedKey[98]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_98_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_98_n29), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_98_n28), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_98_n27), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_98_n30) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_98_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n82), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_98_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n87), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_98_n27) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_98_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n82), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_98_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n87), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_98_n28) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_98_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_98_n25), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n71), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_98_n26) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_98_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n58), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_98_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_98_n25) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_98_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n71), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_98_n23), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n58), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_98_n29) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_98_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_98_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_98_n23) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_98_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n58), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_98_n24) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_99_U9 ( .A(
        KeyMux_D0_input[99]), .B(KeyMux_D1_input[99]), .S(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_99_n30), .Z(Red_SelectedKey[99]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_99_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_99_n29), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_99_n28), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_99_n27), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_99_n30) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_99_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n82), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_99_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n87), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_99_n27) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_99_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n82), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_99_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n87), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_99_n28) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_99_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_99_n25), .B(n3), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_99_n26) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_99_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n63), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_99_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_99_n25) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_99_U3 ( .A1(n3), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_99_n23), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n63), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_99_n29) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_99_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_99_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_99_n23) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_99_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n63), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_99_n24) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_100_U9 ( .A(
        KeyMux_D0_input[100]), .B(KeyMux_D1_input[100]), .S(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_100_n30), .Z(
        Red_SelectedKey[100]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_100_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_100_n29), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_100_n28), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_100_n27), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_100_n30) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_100_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n82), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_100_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n87), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_100_n27) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_100_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n82), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_100_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n87), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_100_n28) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_100_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_100_n25), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n69), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_100_n26) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_100_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n63), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_100_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_100_n25) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_100_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n69), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_100_n23), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n63), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_100_n29) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_100_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_100_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_100_n23) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_100_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n63), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_100_n24) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_101_U9 ( .A(
        KeyMux_D0_input[101]), .B(KeyMux_D1_input[101]), .S(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_101_n31), .Z(
        Red_SelectedKey[101]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_101_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_101_n30), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_101_n29), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_101_n28), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_101_n31) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_101_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n82), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_101_n27), .A3(n7), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_101_n28) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_101_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n82), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_101_n27), .A3(n7), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_101_n29) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_101_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_101_n26), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n71), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_101_n27) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_101_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n59), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_101_n25), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_101_n26) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_101_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n71), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_101_n24), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n59), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_101_n30) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_101_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_101_n25), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_101_n24) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_101_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n59), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_101_n25) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_102_U9 ( .A(
        KeyMux_D0_input[102]), .B(KeyMux_D1_input[102]), .S(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_102_n30), .Z(
        Red_SelectedKey[102]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_102_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_102_n29), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_102_n28), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_102_n27), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_102_n30) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_102_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n82), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_102_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n88), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_102_n27) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_102_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n82), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_102_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n88), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_102_n28) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_102_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_102_n25), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n71), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_102_n26) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_102_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n58), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_102_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_102_n25) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_102_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n71), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_102_n23), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n58), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_102_n29) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_102_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_102_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_102_n23) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_102_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n58), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_102_n24) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_103_U9 ( .A(
        KeyMux_D0_input[103]), .B(KeyMux_D1_input[103]), .S(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_103_n30), .Z(
        Red_SelectedKey[103]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_103_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_103_n29), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_103_n28), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_103_n27), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_103_n30) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_103_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n82), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_103_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n88), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_103_n27) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_103_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n82), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_103_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n88), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_103_n28) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_103_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_103_n25), .B(n3), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_103_n26) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_103_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_103_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_103_n25) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_103_U3 ( .A1(n3), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_103_n23), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_103_n29) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_103_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_103_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_103_n23) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_103_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_103_n24) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_104_U9 ( .A(
        KeyMux_D0_input[104]), .B(KeyMux_D1_input[104]), .S(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_104_n31), .Z(
        Red_SelectedKey[104]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_104_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_104_n30), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_104_n29), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_104_n28), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_104_n31) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_104_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n82), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_104_n27), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n85), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_104_n28) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_104_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n82), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_104_n27), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n85), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_104_n29) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_104_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_104_n26), .B(n3), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_104_n27) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_104_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n59), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_104_n25), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_104_n26) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_104_U3 ( .A1(n3), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_104_n24), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n59), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_104_n30) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_104_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_104_n25), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_104_n24) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_104_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n59), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_104_n25) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_105_U9 ( .A(
        KeyMux_D0_input[105]), .B(KeyMux_D1_input[105]), .S(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_105_n30), .Z(
        Red_SelectedKey[105]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_105_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_105_n29), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_105_n28), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_105_n27), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_105_n30) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_105_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n82), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_105_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n88), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_105_n27) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_105_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n82), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_105_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n88), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_105_n28) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_105_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_105_n25), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n70), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_105_n26) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_105_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n58), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_105_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_105_n25) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_105_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n70), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_105_n23), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n58), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_105_n29) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_105_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_105_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_105_n23) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_105_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n58), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_105_n24) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_106_U9 ( .A(
        KeyMux_D0_input[106]), .B(KeyMux_D1_input[106]), .S(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_106_n30), .Z(
        Red_SelectedKey[106]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_106_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_106_n29), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_106_n28), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_106_n27), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_106_n30) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_106_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n82), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_106_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n85), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_106_n27) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_106_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n82), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_106_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n85), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_106_n28) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_106_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_106_n25), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n70), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_106_n26) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_106_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n63), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_106_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_106_n25) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_106_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n70), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_106_n23), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n63), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_106_n29) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_106_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_106_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_106_n23) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_106_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n63), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_106_n24) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_107_U9 ( .A(
        KeyMux_D0_input[107]), .B(KeyMux_D1_input[107]), .S(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_107_n31), .Z(
        Red_SelectedKey[107]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_107_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_107_n30), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_107_n29), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_107_n28), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_107_n31) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_107_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n82), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_107_n27), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n88), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_107_n28) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_107_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n82), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_107_n27), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n88), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_107_n29) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_107_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_107_n26), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n71), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_107_n27) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_107_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n59), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_107_n25), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_107_n26) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_107_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n71), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_107_n24), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n59), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_107_n30) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_107_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_107_n25), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_107_n24) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_107_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n59), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_107_n25) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_108_U9 ( .A(
        KeyMux_D0_input[108]), .B(KeyMux_D1_input[108]), .S(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_108_n30), .Z(
        Red_SelectedKey[108]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_108_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_108_n29), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_108_n28), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_108_n27), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_108_n30) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_108_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n82), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_108_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n88), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_108_n27) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_108_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n82), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_108_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n88), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_108_n28) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_108_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_108_n25), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n70), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_108_n26) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_108_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_108_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_108_n25) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_108_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n70), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_108_n23), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_108_n29) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_108_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_108_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_108_n23) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_108_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_108_n24) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_109_U9 ( .A(
        KeyMux_D0_input[109]), .B(KeyMux_D1_input[109]), .S(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_109_n30), .Z(
        Red_SelectedKey[109]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_109_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_109_n29), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_109_n28), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_109_n27), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_109_n30) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_109_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n82), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_109_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n85), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_109_n27) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_109_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n82), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_109_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n85), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_109_n28) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_109_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_109_n25), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n70), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_109_n26) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_109_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n60), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_109_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_109_n25) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_109_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n70), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_109_n23), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n60), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_109_n29) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_109_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_109_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_109_n23) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_109_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n60), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_109_n24) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_110_U9 ( .A(
        KeyMux_D0_input[110]), .B(KeyMux_D1_input[110]), .S(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_110_n31), .Z(
        Red_SelectedKey[110]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_110_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_110_n30), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_110_n29), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_110_n28), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_110_n31) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_110_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n82), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_110_n27), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n88), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_110_n28) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_110_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n82), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_110_n27), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n88), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_110_n29) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_110_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_110_n26), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n69), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_110_n27) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_110_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n59), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_110_n25), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_110_n26) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_110_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n69), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_110_n24), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n59), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_110_n30) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_110_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_110_n25), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_110_n24) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_110_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n59), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_110_n25) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_111_U9 ( .A(
        KeyMux_D0_input[111]), .B(KeyMux_D1_input[111]), .S(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_111_n30), .Z(
        Red_SelectedKey[111]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_111_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_111_n29), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_111_n28), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_111_n27), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_111_n30) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_111_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n82), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_111_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n85), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_111_n27) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_111_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n82), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_111_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n85), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_111_n28) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_111_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_111_n25), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n69), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_111_n26) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_111_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n60), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_111_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_111_n25) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_111_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n69), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_111_n23), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n60), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_111_n29) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_111_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_111_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_111_n23) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_111_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n60), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_111_n24) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_112_U9 ( .A(Key[64]), .B(
        Key[0]), .S(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_112_n30), .Z(
        SelectedKey[0]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_112_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_112_n29), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_112_n28), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_112_n27), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_112_n30) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_112_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n74), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_112_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n89), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_112_n27) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_112_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n74), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_112_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n89), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_112_n28) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_112_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_112_n25), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n70), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_112_n26) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_112_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n63), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_112_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_112_n25) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_112_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n70), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_112_n23), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n63), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_112_n29) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_112_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_112_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_112_n23) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_112_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n63), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_112_n24) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_113_U9 ( .A(Key[65]), .B(
        Key[1]), .S(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_113_n30), .Z(
        SelectedKey[1]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_113_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_113_n29), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_113_n28), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_113_n27), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_113_n30) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_113_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n73), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_113_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n84), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_113_n27) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_113_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n73), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_113_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n84), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_113_n28) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_113_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_113_n25), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n66), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_113_n26) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_113_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n61), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_113_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_113_n25) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_113_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n66), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_113_n23), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n61), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_113_n29) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_113_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_113_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_113_n23) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_113_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n61), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_113_n24) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_114_U9 ( .A(Key[66]), .B(
        Key[2]), .S(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_114_n30), .Z(
        SelectedKey[2]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_114_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_114_n29), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_114_n28), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_114_n27), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_114_n30) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_114_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n78), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_114_n26), .A3(n7), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_114_n27) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_114_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n78), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_114_n26), .A3(n7), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_114_n28) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_114_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_114_n25), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n66), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_114_n26) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_114_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n63), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_114_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_114_n25) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_114_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n66), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_114_n23), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n63), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_114_n29) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_114_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_114_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_114_n23) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_114_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n63), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_114_n24) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_115_U9 ( .A(Key[67]), .B(
        Key[3]), .S(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_115_n30), .Z(
        SelectedKey[3]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_115_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_115_n29), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_115_n28), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_115_n27), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_115_n30) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_115_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n81), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_115_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n89), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_115_n27) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_115_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n81), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_115_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n89), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_115_n28) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_115_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_115_n25), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n70), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_115_n26) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_115_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_115_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_115_n25) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_115_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n70), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_115_n23), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_115_n29) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_115_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_115_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_115_n23) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_115_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_115_n24) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_116_U9 ( .A(Key[68]), .B(
        Key[4]), .S(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_116_n30), .Z(
        SelectedKey[4]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_116_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_116_n29), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_116_n28), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_116_n27), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_116_n30) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_116_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n77), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_116_n26), .A3(n7), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_116_n27) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_116_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n77), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_116_n26), .A3(n7), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_116_n28) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_116_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_116_n25), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n66), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_116_n26) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_116_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n60), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_116_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_116_n25) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_116_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n66), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_116_n23), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n60), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_116_n29) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_116_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_116_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_116_n23) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_116_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n60), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_116_n24) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_117_U9 ( .A(Key[69]), .B(
        Key[5]), .S(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_117_n30), .Z(
        SelectedKey[5]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_117_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_117_n29), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_117_n28), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_117_n27), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_117_n30) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_117_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n78), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_117_n26), .A3(n7), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_117_n27) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_117_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n78), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_117_n26), .A3(n7), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_117_n28) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_117_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_117_n25), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n66), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_117_n26) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_117_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n60), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_117_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_117_n25) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_117_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n66), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_117_n23), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n60), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_117_n29) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_117_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_117_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_117_n23) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_117_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n60), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_117_n24) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_118_U9 ( .A(Key[70]), .B(
        Key[6]), .S(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_118_n30), .Z(
        SelectedKey[6]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_118_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_118_n29), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_118_n28), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_118_n27), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_118_n30) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_118_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n78), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_118_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n84), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_118_n27) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_118_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n78), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_118_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n84), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_118_n28) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_118_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_118_n25), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n70), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_118_n26) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_118_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n61), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_118_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_118_n25) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_118_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n70), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_118_n23), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n61), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_118_n29) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_118_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_118_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_118_n23) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_118_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n61), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_118_n24) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_119_U9 ( .A(Key[71]), .B(
        Key[7]), .S(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_119_n30), .Z(
        SelectedKey[7]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_119_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_119_n29), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_119_n28), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_119_n27), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_119_n30) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_119_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n77), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_119_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n86), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_119_n27) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_119_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n77), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_119_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n86), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_119_n28) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_119_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_119_n25), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n70), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_119_n26) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_119_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n61), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_119_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_119_n25) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_119_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n70), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_119_n23), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n61), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_119_n29) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_119_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_119_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_119_n23) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_119_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n61), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_119_n24) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_120_U9 ( .A(Key[72]), .B(
        Key[8]), .S(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_120_n30), .Z(
        SelectedKey[8]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_120_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_120_n29), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_120_n28), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_120_n27), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_120_n30) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_120_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n78), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_120_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n85), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_120_n27) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_120_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n78), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_120_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n85), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_120_n28) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_120_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_120_n25), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n70), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_120_n26) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_120_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n61), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_120_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_120_n25) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_120_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n70), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_120_n23), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n61), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_120_n29) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_120_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_120_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_120_n23) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_120_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n61), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_120_n24) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_121_U9 ( .A(Key[73]), .B(
        Key[9]), .S(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_121_n30), .Z(
        SelectedKey[9]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_121_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_121_n29), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_121_n28), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_121_n27), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_121_n30) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_121_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n78), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_121_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n86), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_121_n27) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_121_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n78), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_121_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n86), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_121_n28) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_121_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_121_n25), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n70), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_121_n26) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_121_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n61), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_121_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_121_n25) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_121_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n70), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_121_n23), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n61), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_121_n29) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_121_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_121_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_121_n23) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_121_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n61), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_121_n24) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_122_U9 ( .A(Key[74]), .B(
        Key[10]), .S(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_122_n30), .Z(
        SelectedKey[10]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_122_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_122_n29), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_122_n28), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_122_n27), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_122_n30) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_122_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n78), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_122_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n89), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_122_n27) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_122_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n78), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_122_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n89), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_122_n28) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_122_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_122_n25), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n70), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_122_n26) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_122_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n61), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_122_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_122_n25) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_122_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n70), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_122_n23), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n61), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_122_n29) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_122_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_122_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_122_n23) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_122_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n61), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_122_n24) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_123_U9 ( .A(Key[75]), .B(
        Key[11]), .S(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_123_n30), .Z(
        SelectedKey[11]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_123_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_123_n29), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_123_n28), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_123_n27), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_123_n30) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_123_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n77), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_123_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n83), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_123_n27) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_123_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n77), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_123_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n83), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_123_n28) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_123_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_123_n25), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n70), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_123_n26) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_123_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n61), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_123_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_123_n25) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_123_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n70), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_123_n23), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n61), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_123_n29) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_123_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_123_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_123_n23) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_123_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n61), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_123_n24) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_124_U9 ( .A(Key[76]), .B(
        Key[12]), .S(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_124_n30), .Z(
        SelectedKey[12]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_124_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_124_n29), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_124_n28), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_124_n27), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_124_n30) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_124_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n78), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_124_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n84), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_124_n27) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_124_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n78), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_124_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n84), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_124_n28) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_124_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_124_n25), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n70), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_124_n26) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_124_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n61), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_124_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_124_n25) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_124_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n70), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_124_n23), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n61), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_124_n29) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_124_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_124_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_124_n23) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_124_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n61), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_124_n24) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_125_U9 ( .A(Key[77]), .B(
        Key[13]), .S(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_125_n30), .Z(
        SelectedKey[13]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_125_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_125_n29), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_125_n28), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_125_n27), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_125_n30) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_125_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n78), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_125_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n83), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_125_n27) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_125_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n78), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_125_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n83), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_125_n28) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_125_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_125_n25), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n70), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_125_n26) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_125_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n61), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_125_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_125_n25) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_125_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n70), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_125_n23), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n61), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_125_n29) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_125_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_125_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_125_n23) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_125_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n61), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_125_n24) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_126_U9 ( .A(Key[78]), .B(
        Key[14]), .S(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_126_n30), .Z(
        SelectedKey[14]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_126_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_126_n29), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_126_n28), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_126_n27), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_126_n30) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_126_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n78), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_126_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n86), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_126_n27) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_126_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n78), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_126_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n86), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_126_n28) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_126_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_126_n25), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n70), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_126_n26) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_126_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n61), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_126_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_126_n25) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_126_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n70), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_126_n23), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n61), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_126_n29) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_126_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_126_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_126_n23) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_126_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n61), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_126_n24) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_127_U9 ( .A(Key[79]), .B(
        Key[15]), .S(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_127_n30), .Z(
        SelectedKey[15]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_127_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_127_n29), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_127_n28), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_127_n27), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_127_n30) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_127_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n78), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_127_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n86), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_127_n27) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_127_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n78), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_127_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n86), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_127_n28) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_127_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_127_n25), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n70), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_127_n26) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_127_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n61), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_127_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_127_n25) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_127_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n70), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_127_n23), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n61), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_127_n29) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_127_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_127_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_127_n23) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_127_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n61), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_127_n24) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_128_U9 ( .A(Key[80]), .B(
        Key[16]), .S(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_128_n30), .Z(
        SelectedKey[16]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_128_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_128_n29), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_128_n28), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_128_n27), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_128_n30) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_128_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n78), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_128_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n84), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_128_n27) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_128_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n78), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_128_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n84), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_128_n28) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_128_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_128_n25), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n70), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_128_n26) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_128_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n61), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_128_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_128_n25) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_128_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n70), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_128_n23), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n61), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_128_n29) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_128_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_128_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_128_n23) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_128_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n61), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_128_n24) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_129_U9 ( .A(Key[81]), .B(
        Key[17]), .S(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_129_n30), .Z(
        SelectedKey[17]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_129_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_129_n29), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_129_n28), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_129_n27), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_129_n30) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_129_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n78), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_129_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n85), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_129_n27) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_129_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n78), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_129_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n85), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_129_n28) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_129_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_129_n25), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n70), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_129_n26) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_129_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n61), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_129_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_129_n25) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_129_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n70), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_129_n23), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n61), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_129_n29) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_129_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_129_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_129_n23) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_129_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n61), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_129_n24) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_130_U9 ( .A(Key[82]), .B(
        Key[18]), .S(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_130_n30), .Z(
        SelectedKey[18]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_130_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_130_n29), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_130_n28), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_130_n27), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_130_n30) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_130_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n79), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_130_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n87), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_130_n27) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_130_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n79), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_130_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n87), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_130_n28) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_130_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_130_n25), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n71), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_130_n26) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_130_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n60), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_130_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_130_n25) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_130_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n71), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_130_n23), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n60), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_130_n29) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_130_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_130_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_130_n23) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_130_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n60), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_130_n24) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_131_U9 ( .A(Key[83]), .B(
        Key[19]), .S(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_131_n30), .Z(
        SelectedKey[19]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_131_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_131_n29), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_131_n28), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_131_n27), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_131_n30) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_131_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n79), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_131_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n87), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_131_n27) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_131_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n79), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_131_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n87), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_131_n28) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_131_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_131_n25), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n71), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_131_n26) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_131_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_131_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_131_n25) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_131_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n71), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_131_n23), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_131_n29) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_131_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_131_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_131_n23) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_131_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_131_n24) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_132_U9 ( .A(Key[84]), .B(
        Key[20]), .S(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_132_n30), .Z(
        SelectedKey[20]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_132_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_132_n29), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_132_n28), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_132_n27), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_132_n30) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_132_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n79), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_132_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n87), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_132_n27) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_132_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n79), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_132_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n87), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_132_n28) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_132_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_132_n25), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n71), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_132_n26) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_132_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n60), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_132_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_132_n25) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_132_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n71), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_132_n23), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n60), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_132_n29) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_132_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_132_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_132_n23) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_132_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n60), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_132_n24) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_133_U9 ( .A(Key[85]), .B(
        Key[21]), .S(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_133_n30), .Z(
        SelectedKey[21]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_133_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_133_n29), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_133_n28), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_133_n27), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_133_n30) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_133_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n79), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_133_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n87), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_133_n27) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_133_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n79), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_133_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n87), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_133_n28) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_133_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_133_n25), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n71), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_133_n26) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_133_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_133_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_133_n25) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_133_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n71), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_133_n23), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_133_n29) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_133_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_133_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_133_n23) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_133_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_133_n24) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_134_U9 ( .A(Key[86]), .B(
        Key[22]), .S(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_134_n30), .Z(
        SelectedKey[22]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_134_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_134_n29), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_134_n28), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_134_n27), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_134_n30) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_134_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n79), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_134_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n87), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_134_n27) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_134_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n79), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_134_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n87), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_134_n28) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_134_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_134_n25), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n71), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_134_n26) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_134_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n63), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_134_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_134_n25) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_134_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n71), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_134_n23), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n63), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_134_n29) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_134_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_134_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_134_n23) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_134_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n63), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_134_n24) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_135_U9 ( .A(Key[87]), .B(
        Key[23]), .S(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_135_n30), .Z(
        SelectedKey[23]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_135_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_135_n29), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_135_n28), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_135_n27), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_135_n30) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_135_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n79), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_135_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n87), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_135_n27) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_135_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n79), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_135_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n87), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_135_n28) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_135_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_135_n25), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n71), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_135_n26) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_135_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_135_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_135_n25) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_135_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n71), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_135_n23), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_135_n29) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_135_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_135_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_135_n23) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_135_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_135_n24) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_136_U9 ( .A(Key[88]), .B(
        Key[24]), .S(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_136_n30), .Z(
        SelectedKey[24]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_136_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_136_n29), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_136_n28), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_136_n27), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_136_n30) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_136_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n79), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_136_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n87), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_136_n27) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_136_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n79), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_136_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n87), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_136_n28) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_136_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_136_n25), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n71), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_136_n26) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_136_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n63), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_136_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_136_n25) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_136_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n71), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_136_n23), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n63), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_136_n29) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_136_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_136_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_136_n23) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_136_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n63), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_136_n24) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_137_U9 ( .A(Key[89]), .B(
        Key[25]), .S(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_137_n30), .Z(
        SelectedKey[25]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_137_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_137_n29), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_137_n28), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_137_n27), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_137_n30) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_137_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n79), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_137_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n87), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_137_n27) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_137_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n79), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_137_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n87), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_137_n28) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_137_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_137_n25), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n71), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_137_n26) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_137_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n60), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_137_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_137_n25) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_137_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n71), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_137_n23), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n60), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_137_n29) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_137_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_137_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_137_n23) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_137_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n60), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_137_n24) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_138_U9 ( .A(Key[90]), .B(
        Key[26]), .S(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_138_n30), .Z(
        SelectedKey[26]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_138_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_138_n29), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_138_n28), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_138_n27), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_138_n30) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_138_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n79), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_138_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n87), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_138_n27) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_138_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n79), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_138_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n87), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_138_n28) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_138_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_138_n25), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n71), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_138_n26) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_138_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_138_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_138_n25) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_138_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n71), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_138_n23), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_138_n29) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_138_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_138_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_138_n23) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_138_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_138_n24) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_139_U9 ( .A(Key[91]), .B(
        Key[27]), .S(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_139_n30), .Z(
        SelectedKey[27]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_139_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_139_n29), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_139_n28), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_139_n27), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_139_n30) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_139_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n79), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_139_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n87), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_139_n27) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_139_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n79), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_139_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n87), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_139_n28) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_139_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_139_n25), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n71), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_139_n26) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_139_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n63), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_139_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_139_n25) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_139_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n71), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_139_n23), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n63), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_139_n29) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_139_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_139_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_139_n23) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_139_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n63), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_139_n24) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_140_U9 ( .A(Key[92]), .B(
        Key[28]), .S(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_140_n30), .Z(
        SelectedKey[28]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_140_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_140_n29), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_140_n28), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_140_n27), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_140_n30) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_140_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n79), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_140_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n87), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_140_n27) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_140_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n79), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_140_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n87), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_140_n28) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_140_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_140_n25), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n71), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_140_n26) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_140_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n60), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_140_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_140_n25) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_140_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n71), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_140_n23), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n60), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_140_n29) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_140_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_140_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_140_n23) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_140_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n60), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_140_n24) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_141_U9 ( .A(Key[93]), .B(
        Key[29]), .S(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_141_n30), .Z(
        SelectedKey[29]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_141_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_141_n29), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_141_n28), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_141_n27), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_141_n30) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_141_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n79), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_141_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n87), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_141_n27) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_141_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n79), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_141_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n87), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_141_n28) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_141_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_141_n25), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n71), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_141_n26) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_141_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_141_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_141_n25) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_141_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n71), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_141_n23), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_141_n29) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_141_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_141_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_141_n23) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_141_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_141_n24) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_142_U9 ( .A(Key[94]), .B(
        Key[30]), .S(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_142_n30), .Z(
        SelectedKey[30]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_142_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_142_n29), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_142_n28), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_142_n27), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_142_n30) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_142_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n80), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_142_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n87), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_142_n27) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_142_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n80), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_142_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n87), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_142_n28) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_142_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_142_n25), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n71), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_142_n26) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_142_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_142_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_142_n25) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_142_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n71), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_142_n23), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_142_n29) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_142_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_142_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_142_n23) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_142_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_142_n24) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_143_U9 ( .A(Key[95]), .B(
        Key[31]), .S(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_143_n30), .Z(
        SelectedKey[31]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_143_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_143_n29), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_143_n28), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_143_n27), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_143_n30) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_143_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n80), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_143_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n86), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_143_n27) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_143_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n80), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_143_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n86), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_143_n28) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_143_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_143_n25), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n71), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_143_n26) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_143_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n60), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_143_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_143_n25) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_143_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n71), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_143_n23), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n60), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_143_n29) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_143_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_143_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_143_n23) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_143_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n60), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_143_n24) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_144_U9 ( .A(Key[96]), .B(
        Key[32]), .S(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_144_n30), .Z(
        SelectedKey[32]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_144_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_144_n29), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_144_n28), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_144_n27), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_144_n30) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_144_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n82), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_144_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n88), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_144_n27) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_144_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n82), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_144_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n88), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_144_n28) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_144_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_144_n25), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n69), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_144_n26) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_144_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n58), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_144_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_144_n25) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_144_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n69), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_144_n23), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n58), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_144_n29) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_144_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_144_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_144_n23) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_144_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n58), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_144_n24) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_145_U9 ( .A(Key[97]), .B(
        Key[33]), .S(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_145_n30), .Z(
        SelectedKey[33]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_145_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_145_n29), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_145_n28), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_145_n27), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_145_n30) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_145_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n82), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_145_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n84), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_145_n27) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_145_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n82), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_145_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n84), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_145_n28) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_145_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_145_n25), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n71), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_145_n26) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_145_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n60), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_145_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_145_n25) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_145_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n71), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_145_n23), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n60), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_145_n29) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_145_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_145_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_145_n23) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_145_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n60), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_145_n24) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_146_U9 ( .A(Key[98]), .B(
        Key[34]), .S(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_146_n30), .Z(
        SelectedKey[34]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_146_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_146_n29), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_146_n28), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_146_n27), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_146_n30) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_146_U7 ( .A1(n4), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_146_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n89), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_146_n27) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_146_U6 ( .A1(n4), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_146_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n89), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_146_n28) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_146_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_146_n25), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n72), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_146_n26) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_146_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n61), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_146_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_146_n25) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_146_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n72), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_146_n23), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n61), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_146_n29) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_146_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_146_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_146_n23) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_146_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n61), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_146_n24) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_147_U9 ( .A(Key[99]), .B(
        Key[35]), .S(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_147_n30), .Z(
        SelectedKey[35]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_147_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_147_n29), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_147_n28), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_147_n27), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_147_n30) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_147_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n78), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_147_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n89), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_147_n27) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_147_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n78), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_147_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n89), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_147_n28) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_147_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_147_n25), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n72), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_147_n26) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_147_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n61), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_147_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_147_n25) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_147_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n72), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_147_n23), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n61), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_147_n29) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_147_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_147_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_147_n23) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_147_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n61), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_147_n24) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_148_U9 ( .A(Key[100]), .B(
        Key[36]), .S(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_148_n30), .Z(
        SelectedKey[36]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_148_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_148_n29), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_148_n28), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_148_n27), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_148_n30) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_148_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n79), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_148_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n89), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_148_n27) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_148_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n79), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_148_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n89), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_148_n28) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_148_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_148_n25), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n72), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_148_n26) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_148_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n59), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_148_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_148_n25) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_148_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n72), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_148_n23), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n59), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_148_n29) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_148_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_148_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_148_n23) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_148_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n59), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_148_n24) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_149_U9 ( .A(Key[101]), .B(
        Key[37]), .S(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_149_n30), .Z(
        SelectedKey[37]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_149_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_149_n29), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_149_n28), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_149_n27), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_149_n30) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_149_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n74), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_149_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n89), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_149_n27) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_149_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n74), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_149_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n89), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_149_n28) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_149_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_149_n25), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n72), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_149_n26) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_149_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n63), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_149_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_149_n25) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_149_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n72), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_149_n23), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n63), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_149_n29) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_149_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_149_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_149_n23) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_149_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n63), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_149_n24) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_150_U9 ( .A(Key[102]), .B(
        Key[38]), .S(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_150_n30), .Z(
        SelectedKey[38]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_150_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_150_n29), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_150_n28), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_150_n27), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_150_n30) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_150_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n81), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_150_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n89), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_150_n27) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_150_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n81), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_150_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n89), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_150_n28) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_150_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_150_n25), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n72), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_150_n26) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_150_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n60), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_150_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_150_n25) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_150_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n72), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_150_n23), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n60), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_150_n29) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_150_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_150_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_150_n23) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_150_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n60), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_150_n24) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_151_U9 ( .A(Key[103]), .B(
        Key[39]), .S(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_151_n30), .Z(
        SelectedKey[39]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_151_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_151_n29), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_151_n28), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_151_n27), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_151_n30) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_151_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n73), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_151_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n89), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_151_n27) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_151_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n73), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_151_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n89), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_151_n28) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_151_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_151_n25), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n72), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_151_n26) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_151_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n61), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_151_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_151_n25) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_151_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n72), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_151_n23), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n61), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_151_n29) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_151_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_151_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_151_n23) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_151_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n61), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_151_n24) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_152_U9 ( .A(Key[104]), .B(
        Key[40]), .S(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_152_n30), .Z(
        SelectedKey[40]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_152_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_152_n29), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_152_n28), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_152_n27), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_152_n30) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_152_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n73), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_152_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n89), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_152_n27) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_152_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n73), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_152_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n89), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_152_n28) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_152_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_152_n25), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n72), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_152_n26) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_152_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_152_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_152_n25) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_152_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n72), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_152_n23), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_152_n29) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_152_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_152_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_152_n23) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_152_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_152_n24) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_153_U9 ( .A(Key[105]), .B(
        Key[41]), .S(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_153_n31), .Z(
        SelectedKey[41]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_153_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_153_n30), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_153_n29), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_153_n28), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_153_n31) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_153_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n75), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_153_n27), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n89), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_153_n28) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_153_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n75), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_153_n27), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n89), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_153_n29) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_153_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_153_n26), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n72), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_153_n27) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_153_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n59), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_153_n25), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_153_n26) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_153_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n72), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_153_n24), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n59), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_153_n30) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_153_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_153_n25), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_153_n24) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_153_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n59), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_153_n25) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_154_U9 ( .A(Key[106]), .B(
        Key[42]), .S(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_154_n31), .Z(
        SelectedKey[42]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_154_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_154_n30), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_154_n29), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_154_n28), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_154_n31) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_154_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n74), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_154_n27), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n89), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_154_n28) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_154_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n74), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_154_n27), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n89), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_154_n29) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_154_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_154_n26), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n72), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_154_n27) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_154_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n59), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_154_n25), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_154_n26) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_154_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n72), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_154_n24), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n59), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_154_n30) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_154_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_154_n25), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_154_n24) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_154_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n59), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_154_n25) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_155_U9 ( .A(Key[107]), .B(
        Key[43]), .S(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_155_n30), .Z(
        SelectedKey[43]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_155_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_155_n29), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_155_n28), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_155_n27), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_155_n30) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_155_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n82), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_155_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n89), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_155_n27) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_155_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n82), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_155_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n89), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_155_n28) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_155_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_155_n25), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n72), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_155_n26) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_155_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n60), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_155_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_155_n25) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_155_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n72), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_155_n23), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n60), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_155_n29) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_155_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_155_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_155_n23) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_155_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n60), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_155_n24) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_156_U9 ( .A(Key[108]), .B(
        Key[44]), .S(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_156_n30), .Z(
        SelectedKey[44]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_156_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_156_n29), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_156_n28), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_156_n27), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_156_n30) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_156_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n80), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_156_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n89), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_156_n27) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_156_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n80), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_156_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n89), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_156_n28) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_156_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_156_n25), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n72), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_156_n26) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_156_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_156_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_156_n25) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_156_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n72), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_156_n23), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_156_n29) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_156_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_156_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_156_n23) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_156_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_156_n24) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_157_U9 ( .A(Key[109]), .B(
        Key[45]), .S(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_157_n30), .Z(
        SelectedKey[45]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_157_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_157_n29), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_157_n28), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_157_n27), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_157_n30) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_157_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n77), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_157_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n89), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_157_n27) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_157_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n77), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_157_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n89), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_157_n28) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_157_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_157_n25), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n72), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_157_n26) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_157_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_157_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_157_n25) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_157_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n72), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_157_n23), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_157_n29) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_157_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_157_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_157_n23) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_157_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_157_n24) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_158_U9 ( .A(Key[110]), .B(
        Key[46]), .S(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_158_n30), .Z(
        SelectedKey[46]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_158_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_158_n29), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_158_n28), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_158_n27), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_158_n30) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_158_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n73), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_158_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n86), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_158_n27) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_158_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n73), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_158_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n86), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_158_n28) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_158_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_158_n25), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n72), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_158_n26) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_158_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(n5), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_158_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_158_n25) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_158_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n72), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_158_n23), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(n5), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_158_n29) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_158_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_158_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_158_n23) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_158_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(n5), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_158_n24) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_159_U9 ( .A(Key[111]), .B(
        Key[47]), .S(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_159_n30), .Z(
        SelectedKey[47]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_159_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_159_n29), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_159_n28), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_159_n27), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_159_n30) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_159_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n80), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_159_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n87), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_159_n27) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_159_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n80), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_159_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n87), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_159_n28) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_159_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_159_n25), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n72), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_159_n26) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_159_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(n5), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_159_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_159_n25) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_159_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n72), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_159_n23), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(n5), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_159_n29) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_159_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_159_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_159_n23) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_159_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(n5), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_159_n24) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_160_U9 ( .A(Key[112]), .B(
        Key[48]), .S(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_160_n30), .Z(
        SelectedKey[48]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_160_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_160_n29), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_160_n28), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_160_n27), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_160_n30) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_160_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n73), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_160_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n83), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_160_n27) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_160_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n73), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_160_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n83), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_160_n28) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_160_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_160_n25), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n72), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_160_n26) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_160_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(n5), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_160_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_160_n25) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_160_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n72), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_160_n23), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(n5), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_160_n29) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_160_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_160_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_160_n23) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_160_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(n5), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_160_n24) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_161_U9 ( .A(Key[113]), .B(
        Key[49]), .S(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_161_n30), .Z(
        SelectedKey[49]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_161_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_161_n29), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_161_n28), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_161_n27), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_161_n30) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_161_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n74), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_161_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n83), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_161_n27) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_161_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n74), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_161_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n83), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_161_n28) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_161_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_161_n25), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n72), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_161_n26) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_161_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_161_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_161_n25) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_161_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n72), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_161_n23), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_161_n29) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_161_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_161_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_161_n23) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_161_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_161_n24) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_162_U9 ( .A(Key[114]), .B(
        Key[50]), .S(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_162_n30), .Z(
        SelectedKey[50]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_162_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_162_n29), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_162_n28), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_162_n27), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_162_n30) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_162_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n81), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_162_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n83), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_162_n27) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_162_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n81), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_162_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n83), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_162_n28) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_162_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_162_n25), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n72), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_162_n26) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_162_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n63), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_162_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_162_n25) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_162_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n72), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_162_n23), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n63), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_162_n29) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_162_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_162_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_162_n23) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_162_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n63), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_162_n24) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_163_U9 ( .A(Key[115]), .B(
        Key[51]), .S(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_163_n30), .Z(
        SelectedKey[51]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_163_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_163_n29), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_163_n28), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_163_n27), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_163_n30) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_163_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n81), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_163_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n83), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_163_n27) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_163_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n81), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_163_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n83), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_163_n28) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_163_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_163_n25), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n72), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_163_n26) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_163_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_163_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_163_n25) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_163_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n72), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_163_n23), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_163_n29) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_163_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_163_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_163_n23) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_163_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_163_n24) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_164_U9 ( .A(Key[116]), .B(
        Key[52]), .S(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_164_n30), .Z(
        SelectedKey[52]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_164_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_164_n29), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_164_n28), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_164_n27), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_164_n30) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_164_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n81), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_164_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n83), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_164_n27) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_164_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n81), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_164_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n83), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_164_n28) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_164_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_164_n25), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n72), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_164_n26) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_164_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_164_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_164_n25) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_164_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n72), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_164_n23), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_164_n29) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_164_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_164_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_164_n23) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_164_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_164_n24) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_165_U9 ( .A(Key[117]), .B(
        Key[53]), .S(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_165_n30), .Z(
        SelectedKey[53]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_165_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_165_n29), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_165_n28), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_165_n27), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_165_n30) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_165_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n74), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_165_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n83), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_165_n27) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_165_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n74), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_165_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n83), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_165_n28) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_165_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_165_n25), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n72), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_165_n26) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_165_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_165_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_165_n25) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_165_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n72), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_165_n23), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_165_n29) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_165_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_165_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_165_n23) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_165_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_165_n24) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_166_U9 ( .A(Key[118]), .B(
        Key[54]), .S(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_166_n31), .Z(
        SelectedKey[54]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_166_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_166_n30), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_166_n29), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_166_n28), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_166_n31) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_166_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n78), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_166_n27), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n86), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_166_n28) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_166_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n78), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_166_n27), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n86), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_166_n29) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_166_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_166_n26), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n68), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_166_n27) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_166_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n59), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_166_n25), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_166_n26) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_166_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n68), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_166_n24), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n59), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_166_n30) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_166_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_166_n25), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_166_n24) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_166_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n59), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_166_n25) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_167_U9 ( .A(Key[119]), .B(
        Key[55]), .S(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_167_n30), .Z(
        SelectedKey[55]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_167_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_167_n29), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_167_n28), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_167_n27), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_167_n30) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_167_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n77), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_167_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n87), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_167_n27) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_167_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n77), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_167_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n87), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_167_n28) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_167_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_167_n25), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n68), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_167_n26) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_167_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_167_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_167_n25) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_167_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n68), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_167_n23), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_167_n29) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_167_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_167_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_167_n23) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_167_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_167_n24) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_168_U9 ( .A(Key[120]), .B(
        Key[56]), .S(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_168_n30), .Z(
        SelectedKey[56]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_168_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_168_n29), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_168_n28), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_168_n27), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_168_n30) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_168_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n73), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_168_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n86), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_168_n27) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_168_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n73), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_168_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n86), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_168_n28) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_168_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_168_n25), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n68), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_168_n26) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_168_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n58), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_168_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_168_n25) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_168_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n68), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_168_n23), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n58), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_168_n29) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_168_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_168_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_168_n23) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_168_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n58), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_168_n24) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_169_U9 ( .A(Key[121]), .B(
        Key[57]), .S(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_169_n30), .Z(
        SelectedKey[57]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_169_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_169_n29), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_169_n28), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_169_n27), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_169_n30) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_169_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n73), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_169_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n87), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_169_n27) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_169_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n73), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_169_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n87), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_169_n28) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_169_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_169_n25), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n68), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_169_n26) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_169_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n63), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_169_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_169_n25) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_169_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n68), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_169_n23), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n63), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_169_n29) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_169_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_169_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_169_n23) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_169_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n63), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_169_n24) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_170_U9 ( .A(Key[122]), .B(
        Key[58]), .S(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_170_n30), .Z(
        SelectedKey[58]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_170_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_170_n29), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_170_n28), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_170_n27), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_170_n30) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_170_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n74), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_170_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n84), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_170_n27) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_170_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n74), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_170_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n84), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_170_n28) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_170_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_170_n25), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n68), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_170_n26) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_170_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_170_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_170_n25) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_170_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n68), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_170_n23), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_170_n29) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_170_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_170_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_170_n23) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_170_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_170_n24) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_171_U9 ( .A(Key[123]), .B(
        Key[59]), .S(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_171_n30), .Z(
        SelectedKey[59]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_171_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_171_n29), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_171_n28), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_171_n27), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_171_n30) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_171_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n74), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_171_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n87), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_171_n27) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_171_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n74), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_171_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n87), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_171_n28) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_171_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_171_n25), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n68), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_171_n26) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_171_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_171_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_171_n25) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_171_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n68), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_171_n23), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_171_n29) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_171_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_171_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_171_n23) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_171_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_171_n24) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_172_U9 ( .A(Key[124]), .B(
        Key[60]), .S(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_172_n30), .Z(
        SelectedKey[60]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_172_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_172_n29), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_172_n28), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_172_n27), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_172_n30) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_172_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n73), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_172_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n86), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_172_n27) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_172_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n73), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_172_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n86), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_172_n28) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_172_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_172_n25), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n72), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_172_n26) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_172_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_172_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_172_n25) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_172_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n72), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_172_n23), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_172_n29) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_172_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_172_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_172_n23) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_172_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_172_n24) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_173_U9 ( .A(Key[125]), .B(
        Key[61]), .S(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_173_n30), .Z(
        SelectedKey[61]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_173_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_173_n29), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_173_n28), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_173_n27), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_173_n30) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_173_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n73), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_173_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n87), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_173_n27) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_173_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n73), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_173_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n87), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_173_n28) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_173_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_173_n25), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n72), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_173_n26) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_173_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_173_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_173_n25) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_173_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n72), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_173_n23), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_173_n29) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_173_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_173_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_173_n23) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_173_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_173_n24) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_174_U9 ( .A(Key[126]), .B(
        Key[62]), .S(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_174_n30), .Z(
        SelectedKey[62]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_174_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_174_n29), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_174_n28), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_174_n27), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_174_n30) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_174_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n75), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_174_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n86), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_174_n27) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_174_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n75), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_174_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n86), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_174_n28) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_174_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_174_n25), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n72), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_174_n26) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_174_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_174_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_174_n25) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_174_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n72), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_174_n23), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_174_n29) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_174_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_174_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_174_n23) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_174_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_174_n24) );
  MUX2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_175_U9 ( .A(Key[127]), .B(
        Key[63]), .S(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_175_n30), .Z(
        SelectedKey[63]) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_175_U8 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_175_n29), .B2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_175_n28), .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_175_n27), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_175_n30) );
  NAND3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_175_U7 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n81), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_175_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n87), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_175_n27) );
  NOR3_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_175_U6 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n81), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_175_n26), .A3(
        K0K1_KeyMUX_And_Red_KeyMUX_n87), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_175_n28) );
  XNOR2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_175_U5 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_175_n25), .B(
        K0K1_KeyMUX_And_Red_KeyMUX_n72), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_175_n26) );
  OAI21_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_175_U4 ( .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .A(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_175_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_175_n25) );
  OAI22_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_175_U3 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n72), .A2(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_175_n23), .B1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .B2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_175_n29) );
  INV_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_175_U2 ( .A(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_175_n24), .ZN(
        K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_175_n23) );
  NAND2_X1 K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_175_U1 ( .A1(
        K0K1_KeyMUX_And_Red_KeyMUX_n64), .A2(K0K1_KeyMUX_And_Red_KeyMUX_n62), 
        .ZN(K0K1_KeyMUX_And_Red_KeyMUX_MUX2to1Inst_175_n24) );
  XNOR2_X1 Red_K0Inst_LFInst_0_LFInst_0_U2 ( .A(
        Red_K0Inst_LFInst_0_LFInst_0_n3), .B(Key[66]), .ZN(KeyMux_D0_input[0])
         );
  XNOR2_X1 Red_K0Inst_LFInst_0_LFInst_0_U1 ( .A(Key[64]), .B(Key[65]), .ZN(
        Red_K0Inst_LFInst_0_LFInst_0_n3) );
  XNOR2_X1 Red_K0Inst_LFInst_0_LFInst_1_U2 ( .A(
        Red_K0Inst_LFInst_0_LFInst_1_n3), .B(Key[67]), .ZN(KeyMux_D0_input[1])
         );
  XNOR2_X1 Red_K0Inst_LFInst_0_LFInst_1_U1 ( .A(Key[64]), .B(Key[65]), .ZN(
        Red_K0Inst_LFInst_0_LFInst_1_n3) );
  XOR2_X1 Red_K0Inst_LFInst_0_LFInst_2_U1 ( .A(Key[64]), .B(Key[66]), .Z(
        KeyMux_D0_input[2]) );
  XOR2_X1 Red_K0Inst_LFInst_0_LFInst_3_U1 ( .A(Key[64]), .B(Key[67]), .Z(
        KeyMux_D0_input[3]) );
  XOR2_X1 Red_K0Inst_LFInst_0_LFInst_4_U1 ( .A(Key[65]), .B(Key[66]), .Z(
        KeyMux_D0_input[4]) );
  XOR2_X1 Red_K0Inst_LFInst_0_LFInst_5_U1 ( .A(Key[65]), .B(Key[67]), .Z(
        KeyMux_D0_input[5]) );
  XOR2_X1 Red_K0Inst_LFInst_0_LFInst_6_U1 ( .A(Key[66]), .B(Key[67]), .Z(
        KeyMux_D0_input[6]) );
  XNOR2_X1 Red_K0Inst_LFInst_1_LFInst_0_U2 ( .A(
        Red_K0Inst_LFInst_1_LFInst_0_n3), .B(Key[70]), .ZN(KeyMux_D0_input[7])
         );
  XNOR2_X1 Red_K0Inst_LFInst_1_LFInst_0_U1 ( .A(Key[68]), .B(Key[69]), .ZN(
        Red_K0Inst_LFInst_1_LFInst_0_n3) );
  XNOR2_X1 Red_K0Inst_LFInst_1_LFInst_1_U2 ( .A(
        Red_K0Inst_LFInst_1_LFInst_1_n3), .B(Key[71]), .ZN(KeyMux_D0_input[8])
         );
  XNOR2_X1 Red_K0Inst_LFInst_1_LFInst_1_U1 ( .A(Key[68]), .B(Key[69]), .ZN(
        Red_K0Inst_LFInst_1_LFInst_1_n3) );
  XOR2_X1 Red_K0Inst_LFInst_1_LFInst_2_U1 ( .A(Key[68]), .B(Key[70]), .Z(
        KeyMux_D0_input[9]) );
  XOR2_X1 Red_K0Inst_LFInst_1_LFInst_3_U1 ( .A(Key[68]), .B(Key[71]), .Z(
        KeyMux_D0_input[10]) );
  XOR2_X1 Red_K0Inst_LFInst_1_LFInst_4_U1 ( .A(Key[69]), .B(Key[70]), .Z(
        KeyMux_D0_input[11]) );
  XOR2_X1 Red_K0Inst_LFInst_1_LFInst_5_U1 ( .A(Key[69]), .B(Key[71]), .Z(
        KeyMux_D0_input[12]) );
  XOR2_X1 Red_K0Inst_LFInst_1_LFInst_6_U1 ( .A(Key[70]), .B(Key[71]), .Z(
        KeyMux_D0_input[13]) );
  XNOR2_X1 Red_K0Inst_LFInst_2_LFInst_0_U2 ( .A(
        Red_K0Inst_LFInst_2_LFInst_0_n3), .B(Key[74]), .ZN(KeyMux_D0_input[14]) );
  XNOR2_X1 Red_K0Inst_LFInst_2_LFInst_0_U1 ( .A(Key[72]), .B(Key[73]), .ZN(
        Red_K0Inst_LFInst_2_LFInst_0_n3) );
  XNOR2_X1 Red_K0Inst_LFInst_2_LFInst_1_U2 ( .A(
        Red_K0Inst_LFInst_2_LFInst_1_n3), .B(Key[75]), .ZN(KeyMux_D0_input[15]) );
  XNOR2_X1 Red_K0Inst_LFInst_2_LFInst_1_U1 ( .A(Key[72]), .B(Key[73]), .ZN(
        Red_K0Inst_LFInst_2_LFInst_1_n3) );
  XOR2_X1 Red_K0Inst_LFInst_2_LFInst_2_U1 ( .A(Key[72]), .B(Key[74]), .Z(
        KeyMux_D0_input[16]) );
  XOR2_X1 Red_K0Inst_LFInst_2_LFInst_3_U1 ( .A(Key[72]), .B(Key[75]), .Z(
        KeyMux_D0_input[17]) );
  XOR2_X1 Red_K0Inst_LFInst_2_LFInst_4_U1 ( .A(Key[73]), .B(Key[74]), .Z(
        KeyMux_D0_input[18]) );
  XOR2_X1 Red_K0Inst_LFInst_2_LFInst_5_U1 ( .A(Key[73]), .B(Key[75]), .Z(
        KeyMux_D0_input[19]) );
  XOR2_X1 Red_K0Inst_LFInst_2_LFInst_6_U1 ( .A(Key[74]), .B(Key[75]), .Z(
        KeyMux_D0_input[20]) );
  XNOR2_X1 Red_K0Inst_LFInst_3_LFInst_0_U2 ( .A(
        Red_K0Inst_LFInst_3_LFInst_0_n3), .B(Key[78]), .ZN(KeyMux_D0_input[21]) );
  XNOR2_X1 Red_K0Inst_LFInst_3_LFInst_0_U1 ( .A(Key[76]), .B(Key[77]), .ZN(
        Red_K0Inst_LFInst_3_LFInst_0_n3) );
  XNOR2_X1 Red_K0Inst_LFInst_3_LFInst_1_U2 ( .A(
        Red_K0Inst_LFInst_3_LFInst_1_n3), .B(Key[79]), .ZN(KeyMux_D0_input[22]) );
  XNOR2_X1 Red_K0Inst_LFInst_3_LFInst_1_U1 ( .A(Key[76]), .B(Key[77]), .ZN(
        Red_K0Inst_LFInst_3_LFInst_1_n3) );
  XOR2_X1 Red_K0Inst_LFInst_3_LFInst_2_U1 ( .A(Key[76]), .B(Key[78]), .Z(
        KeyMux_D0_input[23]) );
  XOR2_X1 Red_K0Inst_LFInst_3_LFInst_3_U1 ( .A(Key[76]), .B(Key[79]), .Z(
        KeyMux_D0_input[24]) );
  XOR2_X1 Red_K0Inst_LFInst_3_LFInst_4_U1 ( .A(Key[77]), .B(Key[78]), .Z(
        KeyMux_D0_input[25]) );
  XOR2_X1 Red_K0Inst_LFInst_3_LFInst_5_U1 ( .A(Key[77]), .B(Key[79]), .Z(
        KeyMux_D0_input[26]) );
  XOR2_X1 Red_K0Inst_LFInst_3_LFInst_6_U1 ( .A(Key[78]), .B(Key[79]), .Z(
        KeyMux_D0_input[27]) );
  XNOR2_X1 Red_K0Inst_LFInst_4_LFInst_0_U2 ( .A(
        Red_K0Inst_LFInst_4_LFInst_0_n3), .B(Key[82]), .ZN(KeyMux_D0_input[28]) );
  XNOR2_X1 Red_K0Inst_LFInst_4_LFInst_0_U1 ( .A(Key[80]), .B(Key[81]), .ZN(
        Red_K0Inst_LFInst_4_LFInst_0_n3) );
  XNOR2_X1 Red_K0Inst_LFInst_4_LFInst_1_U2 ( .A(
        Red_K0Inst_LFInst_4_LFInst_1_n3), .B(Key[83]), .ZN(KeyMux_D0_input[29]) );
  XNOR2_X1 Red_K0Inst_LFInst_4_LFInst_1_U1 ( .A(Key[80]), .B(Key[81]), .ZN(
        Red_K0Inst_LFInst_4_LFInst_1_n3) );
  XOR2_X1 Red_K0Inst_LFInst_4_LFInst_2_U1 ( .A(Key[80]), .B(Key[82]), .Z(
        KeyMux_D0_input[30]) );
  XOR2_X1 Red_K0Inst_LFInst_4_LFInst_3_U1 ( .A(Key[80]), .B(Key[83]), .Z(
        KeyMux_D0_input[31]) );
  XOR2_X1 Red_K0Inst_LFInst_4_LFInst_4_U1 ( .A(Key[81]), .B(Key[82]), .Z(
        KeyMux_D0_input[32]) );
  XOR2_X1 Red_K0Inst_LFInst_4_LFInst_5_U1 ( .A(Key[81]), .B(Key[83]), .Z(
        KeyMux_D0_input[33]) );
  XOR2_X1 Red_K0Inst_LFInst_4_LFInst_6_U1 ( .A(Key[82]), .B(Key[83]), .Z(
        KeyMux_D0_input[34]) );
  XNOR2_X1 Red_K0Inst_LFInst_5_LFInst_0_U2 ( .A(
        Red_K0Inst_LFInst_5_LFInst_0_n3), .B(Key[86]), .ZN(KeyMux_D0_input[35]) );
  XNOR2_X1 Red_K0Inst_LFInst_5_LFInst_0_U1 ( .A(Key[84]), .B(Key[85]), .ZN(
        Red_K0Inst_LFInst_5_LFInst_0_n3) );
  XNOR2_X1 Red_K0Inst_LFInst_5_LFInst_1_U2 ( .A(
        Red_K0Inst_LFInst_5_LFInst_1_n3), .B(Key[87]), .ZN(KeyMux_D0_input[36]) );
  XNOR2_X1 Red_K0Inst_LFInst_5_LFInst_1_U1 ( .A(Key[84]), .B(Key[85]), .ZN(
        Red_K0Inst_LFInst_5_LFInst_1_n3) );
  XOR2_X1 Red_K0Inst_LFInst_5_LFInst_2_U1 ( .A(Key[84]), .B(Key[86]), .Z(
        KeyMux_D0_input[37]) );
  XOR2_X1 Red_K0Inst_LFInst_5_LFInst_3_U1 ( .A(Key[84]), .B(Key[87]), .Z(
        KeyMux_D0_input[38]) );
  XOR2_X1 Red_K0Inst_LFInst_5_LFInst_4_U1 ( .A(Key[85]), .B(Key[86]), .Z(
        KeyMux_D0_input[39]) );
  XOR2_X1 Red_K0Inst_LFInst_5_LFInst_5_U1 ( .A(Key[85]), .B(Key[87]), .Z(
        KeyMux_D0_input[40]) );
  XOR2_X1 Red_K0Inst_LFInst_5_LFInst_6_U1 ( .A(Key[86]), .B(Key[87]), .Z(
        KeyMux_D0_input[41]) );
  XNOR2_X1 Red_K0Inst_LFInst_6_LFInst_0_U2 ( .A(
        Red_K0Inst_LFInst_6_LFInst_0_n3), .B(Key[90]), .ZN(KeyMux_D0_input[42]) );
  XNOR2_X1 Red_K0Inst_LFInst_6_LFInst_0_U1 ( .A(Key[88]), .B(Key[89]), .ZN(
        Red_K0Inst_LFInst_6_LFInst_0_n3) );
  XNOR2_X1 Red_K0Inst_LFInst_6_LFInst_1_U2 ( .A(
        Red_K0Inst_LFInst_6_LFInst_1_n3), .B(Key[91]), .ZN(KeyMux_D0_input[43]) );
  XNOR2_X1 Red_K0Inst_LFInst_6_LFInst_1_U1 ( .A(Key[88]), .B(Key[89]), .ZN(
        Red_K0Inst_LFInst_6_LFInst_1_n3) );
  XOR2_X1 Red_K0Inst_LFInst_6_LFInst_2_U1 ( .A(Key[88]), .B(Key[90]), .Z(
        KeyMux_D0_input[44]) );
  XOR2_X1 Red_K0Inst_LFInst_6_LFInst_3_U1 ( .A(Key[88]), .B(Key[91]), .Z(
        KeyMux_D0_input[45]) );
  XOR2_X1 Red_K0Inst_LFInst_6_LFInst_4_U1 ( .A(Key[89]), .B(Key[90]), .Z(
        KeyMux_D0_input[46]) );
  XOR2_X1 Red_K0Inst_LFInst_6_LFInst_5_U1 ( .A(Key[89]), .B(Key[91]), .Z(
        KeyMux_D0_input[47]) );
  XOR2_X1 Red_K0Inst_LFInst_6_LFInst_6_U1 ( .A(Key[90]), .B(Key[91]), .Z(
        KeyMux_D0_input[48]) );
  XNOR2_X1 Red_K0Inst_LFInst_7_LFInst_0_U2 ( .A(
        Red_K0Inst_LFInst_7_LFInst_0_n3), .B(Key[94]), .ZN(KeyMux_D0_input[49]) );
  XNOR2_X1 Red_K0Inst_LFInst_7_LFInst_0_U1 ( .A(Key[92]), .B(Key[93]), .ZN(
        Red_K0Inst_LFInst_7_LFInst_0_n3) );
  XNOR2_X1 Red_K0Inst_LFInst_7_LFInst_1_U2 ( .A(
        Red_K0Inst_LFInst_7_LFInst_1_n3), .B(Key[95]), .ZN(KeyMux_D0_input[50]) );
  XNOR2_X1 Red_K0Inst_LFInst_7_LFInst_1_U1 ( .A(Key[92]), .B(Key[93]), .ZN(
        Red_K0Inst_LFInst_7_LFInst_1_n3) );
  XOR2_X1 Red_K0Inst_LFInst_7_LFInst_2_U1 ( .A(Key[92]), .B(Key[94]), .Z(
        KeyMux_D0_input[51]) );
  XOR2_X1 Red_K0Inst_LFInst_7_LFInst_3_U1 ( .A(Key[92]), .B(Key[95]), .Z(
        KeyMux_D0_input[52]) );
  XOR2_X1 Red_K0Inst_LFInst_7_LFInst_4_U1 ( .A(Key[93]), .B(Key[94]), .Z(
        KeyMux_D0_input[53]) );
  XOR2_X1 Red_K0Inst_LFInst_7_LFInst_5_U1 ( .A(Key[93]), .B(Key[95]), .Z(
        KeyMux_D0_input[54]) );
  XOR2_X1 Red_K0Inst_LFInst_7_LFInst_6_U1 ( .A(Key[94]), .B(Key[95]), .Z(
        KeyMux_D0_input[55]) );
  XNOR2_X1 Red_K0Inst_LFInst_8_LFInst_0_U2 ( .A(
        Red_K0Inst_LFInst_8_LFInst_0_n3), .B(Key[98]), .ZN(KeyMux_D0_input[56]) );
  XNOR2_X1 Red_K0Inst_LFInst_8_LFInst_0_U1 ( .A(Key[96]), .B(Key[97]), .ZN(
        Red_K0Inst_LFInst_8_LFInst_0_n3) );
  XNOR2_X1 Red_K0Inst_LFInst_8_LFInst_1_U2 ( .A(
        Red_K0Inst_LFInst_8_LFInst_1_n3), .B(Key[99]), .ZN(KeyMux_D0_input[57]) );
  XNOR2_X1 Red_K0Inst_LFInst_8_LFInst_1_U1 ( .A(Key[96]), .B(Key[97]), .ZN(
        Red_K0Inst_LFInst_8_LFInst_1_n3) );
  XOR2_X1 Red_K0Inst_LFInst_8_LFInst_2_U1 ( .A(Key[96]), .B(Key[98]), .Z(
        KeyMux_D0_input[58]) );
  XOR2_X1 Red_K0Inst_LFInst_8_LFInst_3_U1 ( .A(Key[96]), .B(Key[99]), .Z(
        KeyMux_D0_input[59]) );
  XOR2_X1 Red_K0Inst_LFInst_8_LFInst_4_U1 ( .A(Key[97]), .B(Key[98]), .Z(
        KeyMux_D0_input[60]) );
  XOR2_X1 Red_K0Inst_LFInst_8_LFInst_5_U1 ( .A(Key[97]), .B(Key[99]), .Z(
        KeyMux_D0_input[61]) );
  XOR2_X1 Red_K0Inst_LFInst_8_LFInst_6_U1 ( .A(Key[98]), .B(Key[99]), .Z(
        KeyMux_D0_input[62]) );
  XNOR2_X1 Red_K0Inst_LFInst_9_LFInst_0_U2 ( .A(
        Red_K0Inst_LFInst_9_LFInst_0_n3), .B(Key[102]), .ZN(
        KeyMux_D0_input[63]) );
  XNOR2_X1 Red_K0Inst_LFInst_9_LFInst_0_U1 ( .A(Key[100]), .B(Key[101]), .ZN(
        Red_K0Inst_LFInst_9_LFInst_0_n3) );
  XNOR2_X1 Red_K0Inst_LFInst_9_LFInst_1_U2 ( .A(
        Red_K0Inst_LFInst_9_LFInst_1_n3), .B(Key[103]), .ZN(
        KeyMux_D0_input[64]) );
  XNOR2_X1 Red_K0Inst_LFInst_9_LFInst_1_U1 ( .A(Key[100]), .B(Key[101]), .ZN(
        Red_K0Inst_LFInst_9_LFInst_1_n3) );
  XOR2_X1 Red_K0Inst_LFInst_9_LFInst_2_U1 ( .A(Key[100]), .B(Key[102]), .Z(
        KeyMux_D0_input[65]) );
  XOR2_X1 Red_K0Inst_LFInst_9_LFInst_3_U1 ( .A(Key[100]), .B(Key[103]), .Z(
        KeyMux_D0_input[66]) );
  XOR2_X1 Red_K0Inst_LFInst_9_LFInst_4_U1 ( .A(Key[101]), .B(Key[102]), .Z(
        KeyMux_D0_input[67]) );
  XOR2_X1 Red_K0Inst_LFInst_9_LFInst_5_U1 ( .A(Key[101]), .B(Key[103]), .Z(
        KeyMux_D0_input[68]) );
  XOR2_X1 Red_K0Inst_LFInst_9_LFInst_6_U1 ( .A(Key[102]), .B(Key[103]), .Z(
        KeyMux_D0_input[69]) );
  XNOR2_X1 Red_K0Inst_LFInst_10_LFInst_0_U2 ( .A(
        Red_K0Inst_LFInst_10_LFInst_0_n3), .B(Key[106]), .ZN(
        KeyMux_D0_input[70]) );
  XNOR2_X1 Red_K0Inst_LFInst_10_LFInst_0_U1 ( .A(Key[104]), .B(Key[105]), .ZN(
        Red_K0Inst_LFInst_10_LFInst_0_n3) );
  XNOR2_X1 Red_K0Inst_LFInst_10_LFInst_1_U2 ( .A(
        Red_K0Inst_LFInst_10_LFInst_1_n3), .B(Key[107]), .ZN(
        KeyMux_D0_input[71]) );
  XNOR2_X1 Red_K0Inst_LFInst_10_LFInst_1_U1 ( .A(Key[104]), .B(Key[105]), .ZN(
        Red_K0Inst_LFInst_10_LFInst_1_n3) );
  XOR2_X1 Red_K0Inst_LFInst_10_LFInst_2_U1 ( .A(Key[104]), .B(Key[106]), .Z(
        KeyMux_D0_input[72]) );
  XOR2_X1 Red_K0Inst_LFInst_10_LFInst_3_U1 ( .A(Key[104]), .B(Key[107]), .Z(
        KeyMux_D0_input[73]) );
  XOR2_X1 Red_K0Inst_LFInst_10_LFInst_4_U1 ( .A(Key[105]), .B(Key[106]), .Z(
        KeyMux_D0_input[74]) );
  XOR2_X1 Red_K0Inst_LFInst_10_LFInst_5_U1 ( .A(Key[105]), .B(Key[107]), .Z(
        KeyMux_D0_input[75]) );
  XOR2_X1 Red_K0Inst_LFInst_10_LFInst_6_U1 ( .A(Key[106]), .B(Key[107]), .Z(
        KeyMux_D0_input[76]) );
  XNOR2_X1 Red_K0Inst_LFInst_11_LFInst_0_U2 ( .A(
        Red_K0Inst_LFInst_11_LFInst_0_n3), .B(Key[110]), .ZN(
        KeyMux_D0_input[77]) );
  XNOR2_X1 Red_K0Inst_LFInst_11_LFInst_0_U1 ( .A(Key[108]), .B(Key[109]), .ZN(
        Red_K0Inst_LFInst_11_LFInst_0_n3) );
  XNOR2_X1 Red_K0Inst_LFInst_11_LFInst_1_U2 ( .A(
        Red_K0Inst_LFInst_11_LFInst_1_n3), .B(Key[111]), .ZN(
        KeyMux_D0_input[78]) );
  XNOR2_X1 Red_K0Inst_LFInst_11_LFInst_1_U1 ( .A(Key[108]), .B(Key[109]), .ZN(
        Red_K0Inst_LFInst_11_LFInst_1_n3) );
  XOR2_X1 Red_K0Inst_LFInst_11_LFInst_2_U1 ( .A(Key[108]), .B(Key[110]), .Z(
        KeyMux_D0_input[79]) );
  XOR2_X1 Red_K0Inst_LFInst_11_LFInst_3_U1 ( .A(Key[108]), .B(Key[111]), .Z(
        KeyMux_D0_input[80]) );
  XOR2_X1 Red_K0Inst_LFInst_11_LFInst_4_U1 ( .A(Key[109]), .B(Key[110]), .Z(
        KeyMux_D0_input[81]) );
  XOR2_X1 Red_K0Inst_LFInst_11_LFInst_5_U1 ( .A(Key[109]), .B(Key[111]), .Z(
        KeyMux_D0_input[82]) );
  XOR2_X1 Red_K0Inst_LFInst_11_LFInst_6_U1 ( .A(Key[110]), .B(Key[111]), .Z(
        KeyMux_D0_input[83]) );
  XNOR2_X1 Red_K0Inst_LFInst_12_LFInst_0_U2 ( .A(
        Red_K0Inst_LFInst_12_LFInst_0_n3), .B(Key[114]), .ZN(
        KeyMux_D0_input[84]) );
  XNOR2_X1 Red_K0Inst_LFInst_12_LFInst_0_U1 ( .A(Key[112]), .B(Key[113]), .ZN(
        Red_K0Inst_LFInst_12_LFInst_0_n3) );
  XNOR2_X1 Red_K0Inst_LFInst_12_LFInst_1_U2 ( .A(
        Red_K0Inst_LFInst_12_LFInst_1_n3), .B(Key[115]), .ZN(
        KeyMux_D0_input[85]) );
  XNOR2_X1 Red_K0Inst_LFInst_12_LFInst_1_U1 ( .A(Key[112]), .B(Key[113]), .ZN(
        Red_K0Inst_LFInst_12_LFInst_1_n3) );
  XOR2_X1 Red_K0Inst_LFInst_12_LFInst_2_U1 ( .A(Key[112]), .B(Key[114]), .Z(
        KeyMux_D0_input[86]) );
  XOR2_X1 Red_K0Inst_LFInst_12_LFInst_3_U1 ( .A(Key[112]), .B(Key[115]), .Z(
        KeyMux_D0_input[87]) );
  XOR2_X1 Red_K0Inst_LFInst_12_LFInst_4_U1 ( .A(Key[113]), .B(Key[114]), .Z(
        KeyMux_D0_input[88]) );
  XOR2_X1 Red_K0Inst_LFInst_12_LFInst_5_U1 ( .A(Key[113]), .B(Key[115]), .Z(
        KeyMux_D0_input[89]) );
  XOR2_X1 Red_K0Inst_LFInst_12_LFInst_6_U1 ( .A(Key[114]), .B(Key[115]), .Z(
        KeyMux_D0_input[90]) );
  XNOR2_X1 Red_K0Inst_LFInst_13_LFInst_0_U2 ( .A(
        Red_K0Inst_LFInst_13_LFInst_0_n3), .B(Key[118]), .ZN(
        KeyMux_D0_input[91]) );
  XNOR2_X1 Red_K0Inst_LFInst_13_LFInst_0_U1 ( .A(Key[116]), .B(Key[117]), .ZN(
        Red_K0Inst_LFInst_13_LFInst_0_n3) );
  XNOR2_X1 Red_K0Inst_LFInst_13_LFInst_1_U2 ( .A(
        Red_K0Inst_LFInst_13_LFInst_1_n3), .B(Key[119]), .ZN(
        KeyMux_D0_input[92]) );
  XNOR2_X1 Red_K0Inst_LFInst_13_LFInst_1_U1 ( .A(Key[116]), .B(Key[117]), .ZN(
        Red_K0Inst_LFInst_13_LFInst_1_n3) );
  XOR2_X1 Red_K0Inst_LFInst_13_LFInst_2_U1 ( .A(Key[116]), .B(Key[118]), .Z(
        KeyMux_D0_input[93]) );
  XOR2_X1 Red_K0Inst_LFInst_13_LFInst_3_U1 ( .A(Key[116]), .B(Key[119]), .Z(
        KeyMux_D0_input[94]) );
  XOR2_X1 Red_K0Inst_LFInst_13_LFInst_4_U1 ( .A(Key[117]), .B(Key[118]), .Z(
        KeyMux_D0_input[95]) );
  XOR2_X1 Red_K0Inst_LFInst_13_LFInst_5_U1 ( .A(Key[117]), .B(Key[119]), .Z(
        KeyMux_D0_input[96]) );
  XOR2_X1 Red_K0Inst_LFInst_13_LFInst_6_U1 ( .A(Key[118]), .B(Key[119]), .Z(
        KeyMux_D0_input[97]) );
  XNOR2_X1 Red_K0Inst_LFInst_14_LFInst_0_U2 ( .A(
        Red_K0Inst_LFInst_14_LFInst_0_n3), .B(Key[122]), .ZN(
        KeyMux_D0_input[98]) );
  XNOR2_X1 Red_K0Inst_LFInst_14_LFInst_0_U1 ( .A(Key[120]), .B(Key[121]), .ZN(
        Red_K0Inst_LFInst_14_LFInst_0_n3) );
  XNOR2_X1 Red_K0Inst_LFInst_14_LFInst_1_U2 ( .A(
        Red_K0Inst_LFInst_14_LFInst_1_n3), .B(Key[123]), .ZN(
        KeyMux_D0_input[99]) );
  XNOR2_X1 Red_K0Inst_LFInst_14_LFInst_1_U1 ( .A(Key[120]), .B(Key[121]), .ZN(
        Red_K0Inst_LFInst_14_LFInst_1_n3) );
  XOR2_X1 Red_K0Inst_LFInst_14_LFInst_2_U1 ( .A(Key[120]), .B(Key[122]), .Z(
        KeyMux_D0_input[100]) );
  XOR2_X1 Red_K0Inst_LFInst_14_LFInst_3_U1 ( .A(Key[120]), .B(Key[123]), .Z(
        KeyMux_D0_input[101]) );
  XOR2_X1 Red_K0Inst_LFInst_14_LFInst_4_U1 ( .A(Key[121]), .B(Key[122]), .Z(
        KeyMux_D0_input[102]) );
  XOR2_X1 Red_K0Inst_LFInst_14_LFInst_5_U1 ( .A(Key[121]), .B(Key[123]), .Z(
        KeyMux_D0_input[103]) );
  XOR2_X1 Red_K0Inst_LFInst_14_LFInst_6_U1 ( .A(Key[122]), .B(Key[123]), .Z(
        KeyMux_D0_input[104]) );
  XNOR2_X1 Red_K0Inst_LFInst_15_LFInst_0_U2 ( .A(
        Red_K0Inst_LFInst_15_LFInst_0_n3), .B(Key[126]), .ZN(
        KeyMux_D0_input[105]) );
  XNOR2_X1 Red_K0Inst_LFInst_15_LFInst_0_U1 ( .A(Key[124]), .B(Key[125]), .ZN(
        Red_K0Inst_LFInst_15_LFInst_0_n3) );
  XNOR2_X1 Red_K0Inst_LFInst_15_LFInst_1_U2 ( .A(
        Red_K0Inst_LFInst_15_LFInst_1_n3), .B(Key[127]), .ZN(
        KeyMux_D0_input[106]) );
  XNOR2_X1 Red_K0Inst_LFInst_15_LFInst_1_U1 ( .A(Key[124]), .B(Key[125]), .ZN(
        Red_K0Inst_LFInst_15_LFInst_1_n3) );
  XOR2_X1 Red_K0Inst_LFInst_15_LFInst_2_U1 ( .A(Key[124]), .B(Key[126]), .Z(
        KeyMux_D0_input[107]) );
  XOR2_X1 Red_K0Inst_LFInst_15_LFInst_3_U1 ( .A(Key[124]), .B(Key[127]), .Z(
        KeyMux_D0_input[108]) );
  XOR2_X1 Red_K0Inst_LFInst_15_LFInst_4_U1 ( .A(Key[125]), .B(Key[126]), .Z(
        KeyMux_D0_input[109]) );
  XOR2_X1 Red_K0Inst_LFInst_15_LFInst_5_U1 ( .A(Key[125]), .B(Key[127]), .Z(
        KeyMux_D0_input[110]) );
  XOR2_X1 Red_K0Inst_LFInst_15_LFInst_6_U1 ( .A(Key[126]), .B(Key[127]), .Z(
        KeyMux_D0_input[111]) );
  XNOR2_X1 Red_K1Inst_LFInst_0_LFInst_0_U2 ( .A(
        Red_K1Inst_LFInst_0_LFInst_0_n3), .B(Key[2]), .ZN(KeyMux_D1_input[0])
         );
  XNOR2_X1 Red_K1Inst_LFInst_0_LFInst_0_U1 ( .A(Key[0]), .B(Key[1]), .ZN(
        Red_K1Inst_LFInst_0_LFInst_0_n3) );
  XNOR2_X1 Red_K1Inst_LFInst_0_LFInst_1_U2 ( .A(
        Red_K1Inst_LFInst_0_LFInst_1_n3), .B(Key[3]), .ZN(KeyMux_D1_input[1])
         );
  XNOR2_X1 Red_K1Inst_LFInst_0_LFInst_1_U1 ( .A(Key[0]), .B(Key[1]), .ZN(
        Red_K1Inst_LFInst_0_LFInst_1_n3) );
  XOR2_X1 Red_K1Inst_LFInst_0_LFInst_2_U1 ( .A(Key[0]), .B(Key[2]), .Z(
        KeyMux_D1_input[2]) );
  XOR2_X1 Red_K1Inst_LFInst_0_LFInst_3_U1 ( .A(Key[0]), .B(Key[3]), .Z(
        KeyMux_D1_input[3]) );
  XOR2_X1 Red_K1Inst_LFInst_0_LFInst_4_U1 ( .A(Key[1]), .B(Key[2]), .Z(
        KeyMux_D1_input[4]) );
  XOR2_X1 Red_K1Inst_LFInst_0_LFInst_5_U1 ( .A(Key[1]), .B(Key[3]), .Z(
        KeyMux_D1_input[5]) );
  XOR2_X1 Red_K1Inst_LFInst_0_LFInst_6_U1 ( .A(Key[2]), .B(Key[3]), .Z(
        KeyMux_D1_input[6]) );
  XNOR2_X1 Red_K1Inst_LFInst_1_LFInst_0_U2 ( .A(
        Red_K1Inst_LFInst_1_LFInst_0_n3), .B(Key[6]), .ZN(KeyMux_D1_input[7])
         );
  XNOR2_X1 Red_K1Inst_LFInst_1_LFInst_0_U1 ( .A(Key[4]), .B(Key[5]), .ZN(
        Red_K1Inst_LFInst_1_LFInst_0_n3) );
  XNOR2_X1 Red_K1Inst_LFInst_1_LFInst_1_U2 ( .A(
        Red_K1Inst_LFInst_1_LFInst_1_n3), .B(Key[7]), .ZN(KeyMux_D1_input[8])
         );
  XNOR2_X1 Red_K1Inst_LFInst_1_LFInst_1_U1 ( .A(Key[4]), .B(Key[5]), .ZN(
        Red_K1Inst_LFInst_1_LFInst_1_n3) );
  XOR2_X1 Red_K1Inst_LFInst_1_LFInst_2_U1 ( .A(Key[4]), .B(Key[6]), .Z(
        KeyMux_D1_input[9]) );
  XOR2_X1 Red_K1Inst_LFInst_1_LFInst_3_U1 ( .A(Key[4]), .B(Key[7]), .Z(
        KeyMux_D1_input[10]) );
  XOR2_X1 Red_K1Inst_LFInst_1_LFInst_4_U1 ( .A(Key[5]), .B(Key[6]), .Z(
        KeyMux_D1_input[11]) );
  XOR2_X1 Red_K1Inst_LFInst_1_LFInst_5_U1 ( .A(Key[5]), .B(Key[7]), .Z(
        KeyMux_D1_input[12]) );
  XOR2_X1 Red_K1Inst_LFInst_1_LFInst_6_U1 ( .A(Key[6]), .B(Key[7]), .Z(
        KeyMux_D1_input[13]) );
  XNOR2_X1 Red_K1Inst_LFInst_2_LFInst_0_U2 ( .A(
        Red_K1Inst_LFInst_2_LFInst_0_n3), .B(Key[10]), .ZN(KeyMux_D1_input[14]) );
  XNOR2_X1 Red_K1Inst_LFInst_2_LFInst_0_U1 ( .A(Key[8]), .B(Key[9]), .ZN(
        Red_K1Inst_LFInst_2_LFInst_0_n3) );
  XNOR2_X1 Red_K1Inst_LFInst_2_LFInst_1_U2 ( .A(
        Red_K1Inst_LFInst_2_LFInst_1_n3), .B(Key[11]), .ZN(KeyMux_D1_input[15]) );
  XNOR2_X1 Red_K1Inst_LFInst_2_LFInst_1_U1 ( .A(Key[8]), .B(Key[9]), .ZN(
        Red_K1Inst_LFInst_2_LFInst_1_n3) );
  XOR2_X1 Red_K1Inst_LFInst_2_LFInst_2_U1 ( .A(Key[8]), .B(Key[10]), .Z(
        KeyMux_D1_input[16]) );
  XOR2_X1 Red_K1Inst_LFInst_2_LFInst_3_U1 ( .A(Key[8]), .B(Key[11]), .Z(
        KeyMux_D1_input[17]) );
  XOR2_X1 Red_K1Inst_LFInst_2_LFInst_4_U1 ( .A(Key[9]), .B(Key[10]), .Z(
        KeyMux_D1_input[18]) );
  XOR2_X1 Red_K1Inst_LFInst_2_LFInst_5_U1 ( .A(Key[9]), .B(Key[11]), .Z(
        KeyMux_D1_input[19]) );
  XOR2_X1 Red_K1Inst_LFInst_2_LFInst_6_U1 ( .A(Key[10]), .B(Key[11]), .Z(
        KeyMux_D1_input[20]) );
  XNOR2_X1 Red_K1Inst_LFInst_3_LFInst_0_U2 ( .A(
        Red_K1Inst_LFInst_3_LFInst_0_n3), .B(Key[14]), .ZN(KeyMux_D1_input[21]) );
  XNOR2_X1 Red_K1Inst_LFInst_3_LFInst_0_U1 ( .A(Key[12]), .B(Key[13]), .ZN(
        Red_K1Inst_LFInst_3_LFInst_0_n3) );
  XNOR2_X1 Red_K1Inst_LFInst_3_LFInst_1_U2 ( .A(
        Red_K1Inst_LFInst_3_LFInst_1_n3), .B(Key[15]), .ZN(KeyMux_D1_input[22]) );
  XNOR2_X1 Red_K1Inst_LFInst_3_LFInst_1_U1 ( .A(Key[12]), .B(Key[13]), .ZN(
        Red_K1Inst_LFInst_3_LFInst_1_n3) );
  XOR2_X1 Red_K1Inst_LFInst_3_LFInst_2_U1 ( .A(Key[12]), .B(Key[14]), .Z(
        KeyMux_D1_input[23]) );
  XOR2_X1 Red_K1Inst_LFInst_3_LFInst_3_U1 ( .A(Key[12]), .B(Key[15]), .Z(
        KeyMux_D1_input[24]) );
  XOR2_X1 Red_K1Inst_LFInst_3_LFInst_4_U1 ( .A(Key[13]), .B(Key[14]), .Z(
        KeyMux_D1_input[25]) );
  XOR2_X1 Red_K1Inst_LFInst_3_LFInst_5_U1 ( .A(Key[13]), .B(Key[15]), .Z(
        KeyMux_D1_input[26]) );
  XOR2_X1 Red_K1Inst_LFInst_3_LFInst_6_U1 ( .A(Key[14]), .B(Key[15]), .Z(
        KeyMux_D1_input[27]) );
  XNOR2_X1 Red_K1Inst_LFInst_4_LFInst_0_U2 ( .A(
        Red_K1Inst_LFInst_4_LFInst_0_n3), .B(Key[18]), .ZN(KeyMux_D1_input[28]) );
  XNOR2_X1 Red_K1Inst_LFInst_4_LFInst_0_U1 ( .A(Key[16]), .B(Key[17]), .ZN(
        Red_K1Inst_LFInst_4_LFInst_0_n3) );
  XNOR2_X1 Red_K1Inst_LFInst_4_LFInst_1_U2 ( .A(
        Red_K1Inst_LFInst_4_LFInst_1_n3), .B(Key[19]), .ZN(KeyMux_D1_input[29]) );
  XNOR2_X1 Red_K1Inst_LFInst_4_LFInst_1_U1 ( .A(Key[16]), .B(Key[17]), .ZN(
        Red_K1Inst_LFInst_4_LFInst_1_n3) );
  XOR2_X1 Red_K1Inst_LFInst_4_LFInst_2_U1 ( .A(Key[16]), .B(Key[18]), .Z(
        KeyMux_D1_input[30]) );
  XOR2_X1 Red_K1Inst_LFInst_4_LFInst_3_U1 ( .A(Key[16]), .B(Key[19]), .Z(
        KeyMux_D1_input[31]) );
  XOR2_X1 Red_K1Inst_LFInst_4_LFInst_4_U1 ( .A(Key[17]), .B(Key[18]), .Z(
        KeyMux_D1_input[32]) );
  XOR2_X1 Red_K1Inst_LFInst_4_LFInst_5_U1 ( .A(Key[17]), .B(Key[19]), .Z(
        KeyMux_D1_input[33]) );
  XOR2_X1 Red_K1Inst_LFInst_4_LFInst_6_U1 ( .A(Key[18]), .B(Key[19]), .Z(
        KeyMux_D1_input[34]) );
  XNOR2_X1 Red_K1Inst_LFInst_5_LFInst_0_U2 ( .A(
        Red_K1Inst_LFInst_5_LFInst_0_n3), .B(Key[22]), .ZN(KeyMux_D1_input[35]) );
  XNOR2_X1 Red_K1Inst_LFInst_5_LFInst_0_U1 ( .A(Key[20]), .B(Key[21]), .ZN(
        Red_K1Inst_LFInst_5_LFInst_0_n3) );
  XNOR2_X1 Red_K1Inst_LFInst_5_LFInst_1_U2 ( .A(
        Red_K1Inst_LFInst_5_LFInst_1_n3), .B(Key[23]), .ZN(KeyMux_D1_input[36]) );
  XNOR2_X1 Red_K1Inst_LFInst_5_LFInst_1_U1 ( .A(Key[20]), .B(Key[21]), .ZN(
        Red_K1Inst_LFInst_5_LFInst_1_n3) );
  XOR2_X1 Red_K1Inst_LFInst_5_LFInst_2_U1 ( .A(Key[20]), .B(Key[22]), .Z(
        KeyMux_D1_input[37]) );
  XOR2_X1 Red_K1Inst_LFInst_5_LFInst_3_U1 ( .A(Key[20]), .B(Key[23]), .Z(
        KeyMux_D1_input[38]) );
  XOR2_X1 Red_K1Inst_LFInst_5_LFInst_4_U1 ( .A(Key[21]), .B(Key[22]), .Z(
        KeyMux_D1_input[39]) );
  XOR2_X1 Red_K1Inst_LFInst_5_LFInst_5_U1 ( .A(Key[21]), .B(Key[23]), .Z(
        KeyMux_D1_input[40]) );
  XOR2_X1 Red_K1Inst_LFInst_5_LFInst_6_U1 ( .A(Key[22]), .B(Key[23]), .Z(
        KeyMux_D1_input[41]) );
  XNOR2_X1 Red_K1Inst_LFInst_6_LFInst_0_U2 ( .A(
        Red_K1Inst_LFInst_6_LFInst_0_n3), .B(Key[26]), .ZN(KeyMux_D1_input[42]) );
  XNOR2_X1 Red_K1Inst_LFInst_6_LFInst_0_U1 ( .A(Key[24]), .B(Key[25]), .ZN(
        Red_K1Inst_LFInst_6_LFInst_0_n3) );
  XNOR2_X1 Red_K1Inst_LFInst_6_LFInst_1_U2 ( .A(
        Red_K1Inst_LFInst_6_LFInst_1_n3), .B(Key[27]), .ZN(KeyMux_D1_input[43]) );
  XNOR2_X1 Red_K1Inst_LFInst_6_LFInst_1_U1 ( .A(Key[24]), .B(Key[25]), .ZN(
        Red_K1Inst_LFInst_6_LFInst_1_n3) );
  XOR2_X1 Red_K1Inst_LFInst_6_LFInst_2_U1 ( .A(Key[24]), .B(Key[26]), .Z(
        KeyMux_D1_input[44]) );
  XOR2_X1 Red_K1Inst_LFInst_6_LFInst_3_U1 ( .A(Key[24]), .B(Key[27]), .Z(
        KeyMux_D1_input[45]) );
  XOR2_X1 Red_K1Inst_LFInst_6_LFInst_4_U1 ( .A(Key[25]), .B(Key[26]), .Z(
        KeyMux_D1_input[46]) );
  XOR2_X1 Red_K1Inst_LFInst_6_LFInst_5_U1 ( .A(Key[25]), .B(Key[27]), .Z(
        KeyMux_D1_input[47]) );
  XOR2_X1 Red_K1Inst_LFInst_6_LFInst_6_U1 ( .A(Key[26]), .B(Key[27]), .Z(
        KeyMux_D1_input[48]) );
  XNOR2_X1 Red_K1Inst_LFInst_7_LFInst_0_U2 ( .A(
        Red_K1Inst_LFInst_7_LFInst_0_n3), .B(Key[30]), .ZN(KeyMux_D1_input[49]) );
  XNOR2_X1 Red_K1Inst_LFInst_7_LFInst_0_U1 ( .A(Key[28]), .B(Key[29]), .ZN(
        Red_K1Inst_LFInst_7_LFInst_0_n3) );
  XNOR2_X1 Red_K1Inst_LFInst_7_LFInst_1_U2 ( .A(
        Red_K1Inst_LFInst_7_LFInst_1_n3), .B(Key[31]), .ZN(KeyMux_D1_input[50]) );
  XNOR2_X1 Red_K1Inst_LFInst_7_LFInst_1_U1 ( .A(Key[28]), .B(Key[29]), .ZN(
        Red_K1Inst_LFInst_7_LFInst_1_n3) );
  XOR2_X1 Red_K1Inst_LFInst_7_LFInst_2_U1 ( .A(Key[28]), .B(Key[30]), .Z(
        KeyMux_D1_input[51]) );
  XOR2_X1 Red_K1Inst_LFInst_7_LFInst_3_U1 ( .A(Key[28]), .B(Key[31]), .Z(
        KeyMux_D1_input[52]) );
  XOR2_X1 Red_K1Inst_LFInst_7_LFInst_4_U1 ( .A(Key[29]), .B(Key[30]), .Z(
        KeyMux_D1_input[53]) );
  XOR2_X1 Red_K1Inst_LFInst_7_LFInst_5_U1 ( .A(Key[29]), .B(Key[31]), .Z(
        KeyMux_D1_input[54]) );
  XOR2_X1 Red_K1Inst_LFInst_7_LFInst_6_U1 ( .A(Key[30]), .B(Key[31]), .Z(
        KeyMux_D1_input[55]) );
  XNOR2_X1 Red_K1Inst_LFInst_8_LFInst_0_U2 ( .A(
        Red_K1Inst_LFInst_8_LFInst_0_n3), .B(Key[34]), .ZN(KeyMux_D1_input[56]) );
  XNOR2_X1 Red_K1Inst_LFInst_8_LFInst_0_U1 ( .A(Key[32]), .B(Key[33]), .ZN(
        Red_K1Inst_LFInst_8_LFInst_0_n3) );
  XNOR2_X1 Red_K1Inst_LFInst_8_LFInst_1_U2 ( .A(
        Red_K1Inst_LFInst_8_LFInst_1_n3), .B(Key[35]), .ZN(KeyMux_D1_input[57]) );
  XNOR2_X1 Red_K1Inst_LFInst_8_LFInst_1_U1 ( .A(Key[32]), .B(Key[33]), .ZN(
        Red_K1Inst_LFInst_8_LFInst_1_n3) );
  XOR2_X1 Red_K1Inst_LFInst_8_LFInst_2_U1 ( .A(Key[32]), .B(Key[34]), .Z(
        KeyMux_D1_input[58]) );
  XOR2_X1 Red_K1Inst_LFInst_8_LFInst_3_U1 ( .A(Key[32]), .B(Key[35]), .Z(
        KeyMux_D1_input[59]) );
  XOR2_X1 Red_K1Inst_LFInst_8_LFInst_4_U1 ( .A(Key[33]), .B(Key[34]), .Z(
        KeyMux_D1_input[60]) );
  XOR2_X1 Red_K1Inst_LFInst_8_LFInst_5_U1 ( .A(Key[33]), .B(Key[35]), .Z(
        KeyMux_D1_input[61]) );
  XOR2_X1 Red_K1Inst_LFInst_8_LFInst_6_U1 ( .A(Key[34]), .B(Key[35]), .Z(
        KeyMux_D1_input[62]) );
  XNOR2_X1 Red_K1Inst_LFInst_9_LFInst_0_U2 ( .A(
        Red_K1Inst_LFInst_9_LFInst_0_n3), .B(Key[38]), .ZN(KeyMux_D1_input[63]) );
  XNOR2_X1 Red_K1Inst_LFInst_9_LFInst_0_U1 ( .A(Key[36]), .B(Key[37]), .ZN(
        Red_K1Inst_LFInst_9_LFInst_0_n3) );
  XNOR2_X1 Red_K1Inst_LFInst_9_LFInst_1_U2 ( .A(
        Red_K1Inst_LFInst_9_LFInst_1_n3), .B(Key[39]), .ZN(KeyMux_D1_input[64]) );
  XNOR2_X1 Red_K1Inst_LFInst_9_LFInst_1_U1 ( .A(Key[36]), .B(Key[37]), .ZN(
        Red_K1Inst_LFInst_9_LFInst_1_n3) );
  XOR2_X1 Red_K1Inst_LFInst_9_LFInst_2_U1 ( .A(Key[36]), .B(Key[38]), .Z(
        KeyMux_D1_input[65]) );
  XOR2_X1 Red_K1Inst_LFInst_9_LFInst_3_U1 ( .A(Key[36]), .B(Key[39]), .Z(
        KeyMux_D1_input[66]) );
  XOR2_X1 Red_K1Inst_LFInst_9_LFInst_4_U1 ( .A(Key[37]), .B(Key[38]), .Z(
        KeyMux_D1_input[67]) );
  XOR2_X1 Red_K1Inst_LFInst_9_LFInst_5_U1 ( .A(Key[37]), .B(Key[39]), .Z(
        KeyMux_D1_input[68]) );
  XOR2_X1 Red_K1Inst_LFInst_9_LFInst_6_U1 ( .A(Key[38]), .B(Key[39]), .Z(
        KeyMux_D1_input[69]) );
  XNOR2_X1 Red_K1Inst_LFInst_10_LFInst_0_U2 ( .A(
        Red_K1Inst_LFInst_10_LFInst_0_n3), .B(Key[42]), .ZN(
        KeyMux_D1_input[70]) );
  XNOR2_X1 Red_K1Inst_LFInst_10_LFInst_0_U1 ( .A(Key[40]), .B(Key[41]), .ZN(
        Red_K1Inst_LFInst_10_LFInst_0_n3) );
  XNOR2_X1 Red_K1Inst_LFInst_10_LFInst_1_U2 ( .A(
        Red_K1Inst_LFInst_10_LFInst_1_n3), .B(Key[43]), .ZN(
        KeyMux_D1_input[71]) );
  XNOR2_X1 Red_K1Inst_LFInst_10_LFInst_1_U1 ( .A(Key[40]), .B(Key[41]), .ZN(
        Red_K1Inst_LFInst_10_LFInst_1_n3) );
  XOR2_X1 Red_K1Inst_LFInst_10_LFInst_2_U1 ( .A(Key[40]), .B(Key[42]), .Z(
        KeyMux_D1_input[72]) );
  XOR2_X1 Red_K1Inst_LFInst_10_LFInst_3_U1 ( .A(Key[40]), .B(Key[43]), .Z(
        KeyMux_D1_input[73]) );
  XOR2_X1 Red_K1Inst_LFInst_10_LFInst_4_U1 ( .A(Key[41]), .B(Key[42]), .Z(
        KeyMux_D1_input[74]) );
  XOR2_X1 Red_K1Inst_LFInst_10_LFInst_5_U1 ( .A(Key[41]), .B(Key[43]), .Z(
        KeyMux_D1_input[75]) );
  XOR2_X1 Red_K1Inst_LFInst_10_LFInst_6_U1 ( .A(Key[42]), .B(Key[43]), .Z(
        KeyMux_D1_input[76]) );
  XNOR2_X1 Red_K1Inst_LFInst_11_LFInst_0_U2 ( .A(
        Red_K1Inst_LFInst_11_LFInst_0_n3), .B(Key[46]), .ZN(
        KeyMux_D1_input[77]) );
  XNOR2_X1 Red_K1Inst_LFInst_11_LFInst_0_U1 ( .A(Key[44]), .B(Key[45]), .ZN(
        Red_K1Inst_LFInst_11_LFInst_0_n3) );
  XNOR2_X1 Red_K1Inst_LFInst_11_LFInst_1_U2 ( .A(
        Red_K1Inst_LFInst_11_LFInst_1_n3), .B(Key[47]), .ZN(
        KeyMux_D1_input[78]) );
  XNOR2_X1 Red_K1Inst_LFInst_11_LFInst_1_U1 ( .A(Key[44]), .B(Key[45]), .ZN(
        Red_K1Inst_LFInst_11_LFInst_1_n3) );
  XOR2_X1 Red_K1Inst_LFInst_11_LFInst_2_U1 ( .A(Key[44]), .B(Key[46]), .Z(
        KeyMux_D1_input[79]) );
  XOR2_X1 Red_K1Inst_LFInst_11_LFInst_3_U1 ( .A(Key[44]), .B(Key[47]), .Z(
        KeyMux_D1_input[80]) );
  XOR2_X1 Red_K1Inst_LFInst_11_LFInst_4_U1 ( .A(Key[45]), .B(Key[46]), .Z(
        KeyMux_D1_input[81]) );
  XOR2_X1 Red_K1Inst_LFInst_11_LFInst_5_U1 ( .A(Key[45]), .B(Key[47]), .Z(
        KeyMux_D1_input[82]) );
  XOR2_X1 Red_K1Inst_LFInst_11_LFInst_6_U1 ( .A(Key[46]), .B(Key[47]), .Z(
        KeyMux_D1_input[83]) );
  XNOR2_X1 Red_K1Inst_LFInst_12_LFInst_0_U2 ( .A(
        Red_K1Inst_LFInst_12_LFInst_0_n3), .B(Key[50]), .ZN(
        KeyMux_D1_input[84]) );
  XNOR2_X1 Red_K1Inst_LFInst_12_LFInst_0_U1 ( .A(Key[48]), .B(Key[49]), .ZN(
        Red_K1Inst_LFInst_12_LFInst_0_n3) );
  XNOR2_X1 Red_K1Inst_LFInst_12_LFInst_1_U2 ( .A(
        Red_K1Inst_LFInst_12_LFInst_1_n3), .B(Key[51]), .ZN(
        KeyMux_D1_input[85]) );
  XNOR2_X1 Red_K1Inst_LFInst_12_LFInst_1_U1 ( .A(Key[48]), .B(Key[49]), .ZN(
        Red_K1Inst_LFInst_12_LFInst_1_n3) );
  XOR2_X1 Red_K1Inst_LFInst_12_LFInst_2_U1 ( .A(Key[48]), .B(Key[50]), .Z(
        KeyMux_D1_input[86]) );
  XOR2_X1 Red_K1Inst_LFInst_12_LFInst_3_U1 ( .A(Key[48]), .B(Key[51]), .Z(
        KeyMux_D1_input[87]) );
  XOR2_X1 Red_K1Inst_LFInst_12_LFInst_4_U1 ( .A(Key[49]), .B(Key[50]), .Z(
        KeyMux_D1_input[88]) );
  XOR2_X1 Red_K1Inst_LFInst_12_LFInst_5_U1 ( .A(Key[49]), .B(Key[51]), .Z(
        KeyMux_D1_input[89]) );
  XOR2_X1 Red_K1Inst_LFInst_12_LFInst_6_U1 ( .A(Key[50]), .B(Key[51]), .Z(
        KeyMux_D1_input[90]) );
  XNOR2_X1 Red_K1Inst_LFInst_13_LFInst_0_U2 ( .A(
        Red_K1Inst_LFInst_13_LFInst_0_n3), .B(Key[54]), .ZN(
        KeyMux_D1_input[91]) );
  XNOR2_X1 Red_K1Inst_LFInst_13_LFInst_0_U1 ( .A(Key[52]), .B(Key[53]), .ZN(
        Red_K1Inst_LFInst_13_LFInst_0_n3) );
  XNOR2_X1 Red_K1Inst_LFInst_13_LFInst_1_U2 ( .A(
        Red_K1Inst_LFInst_13_LFInst_1_n3), .B(Key[55]), .ZN(
        KeyMux_D1_input[92]) );
  XNOR2_X1 Red_K1Inst_LFInst_13_LFInst_1_U1 ( .A(Key[52]), .B(Key[53]), .ZN(
        Red_K1Inst_LFInst_13_LFInst_1_n3) );
  XOR2_X1 Red_K1Inst_LFInst_13_LFInst_2_U1 ( .A(Key[52]), .B(Key[54]), .Z(
        KeyMux_D1_input[93]) );
  XOR2_X1 Red_K1Inst_LFInst_13_LFInst_3_U1 ( .A(Key[52]), .B(Key[55]), .Z(
        KeyMux_D1_input[94]) );
  XOR2_X1 Red_K1Inst_LFInst_13_LFInst_4_U1 ( .A(Key[53]), .B(Key[54]), .Z(
        KeyMux_D1_input[95]) );
  XOR2_X1 Red_K1Inst_LFInst_13_LFInst_5_U1 ( .A(Key[53]), .B(Key[55]), .Z(
        KeyMux_D1_input[96]) );
  XOR2_X1 Red_K1Inst_LFInst_13_LFInst_6_U1 ( .A(Key[54]), .B(Key[55]), .Z(
        KeyMux_D1_input[97]) );
  XNOR2_X1 Red_K1Inst_LFInst_14_LFInst_0_U2 ( .A(
        Red_K1Inst_LFInst_14_LFInst_0_n3), .B(Key[58]), .ZN(
        KeyMux_D1_input[98]) );
  XNOR2_X1 Red_K1Inst_LFInst_14_LFInst_0_U1 ( .A(Key[56]), .B(Key[57]), .ZN(
        Red_K1Inst_LFInst_14_LFInst_0_n3) );
  XNOR2_X1 Red_K1Inst_LFInst_14_LFInst_1_U2 ( .A(
        Red_K1Inst_LFInst_14_LFInst_1_n3), .B(Key[59]), .ZN(
        KeyMux_D1_input[99]) );
  XNOR2_X1 Red_K1Inst_LFInst_14_LFInst_1_U1 ( .A(Key[56]), .B(Key[57]), .ZN(
        Red_K1Inst_LFInst_14_LFInst_1_n3) );
  XOR2_X1 Red_K1Inst_LFInst_14_LFInst_2_U1 ( .A(Key[56]), .B(Key[58]), .Z(
        KeyMux_D1_input[100]) );
  XOR2_X1 Red_K1Inst_LFInst_14_LFInst_3_U1 ( .A(Key[56]), .B(Key[59]), .Z(
        KeyMux_D1_input[101]) );
  XOR2_X1 Red_K1Inst_LFInst_14_LFInst_4_U1 ( .A(Key[57]), .B(Key[58]), .Z(
        KeyMux_D1_input[102]) );
  XOR2_X1 Red_K1Inst_LFInst_14_LFInst_5_U1 ( .A(Key[57]), .B(Key[59]), .Z(
        KeyMux_D1_input[103]) );
  XOR2_X1 Red_K1Inst_LFInst_14_LFInst_6_U1 ( .A(Key[58]), .B(Key[59]), .Z(
        KeyMux_D1_input[104]) );
  XNOR2_X1 Red_K1Inst_LFInst_15_LFInst_0_U2 ( .A(
        Red_K1Inst_LFInst_15_LFInst_0_n3), .B(Key[62]), .ZN(
        KeyMux_D1_input[105]) );
  XNOR2_X1 Red_K1Inst_LFInst_15_LFInst_0_U1 ( .A(Key[60]), .B(Key[61]), .ZN(
        Red_K1Inst_LFInst_15_LFInst_0_n3) );
  XNOR2_X1 Red_K1Inst_LFInst_15_LFInst_1_U2 ( .A(
        Red_K1Inst_LFInst_15_LFInst_1_n3), .B(Key[63]), .ZN(
        KeyMux_D1_input[106]) );
  XNOR2_X1 Red_K1Inst_LFInst_15_LFInst_1_U1 ( .A(Key[60]), .B(Key[61]), .ZN(
        Red_K1Inst_LFInst_15_LFInst_1_n3) );
  XOR2_X1 Red_K1Inst_LFInst_15_LFInst_2_U1 ( .A(Key[60]), .B(Key[62]), .Z(
        KeyMux_D1_input[107]) );
  XOR2_X1 Red_K1Inst_LFInst_15_LFInst_3_U1 ( .A(Key[60]), .B(Key[63]), .Z(
        KeyMux_D1_input[108]) );
  XOR2_X1 Red_K1Inst_LFInst_15_LFInst_4_U1 ( .A(Key[61]), .B(Key[62]), .Z(
        KeyMux_D1_input[109]) );
  XOR2_X1 Red_K1Inst_LFInst_15_LFInst_5_U1 ( .A(Key[61]), .B(Key[63]), .Z(
        KeyMux_D1_input[110]) );
  XOR2_X1 Red_K1Inst_LFInst_15_LFInst_6_U1 ( .A(Key[62]), .B(Key[63]), .Z(
        KeyMux_D1_input[111]) );
  OR2_X1 FSMMUX_MUXInst_0_U1 ( .A1(FSMReg[0]), .A2(rst), .ZN(FSMF[3]) );
  INV_X1 FSMMUX_MUXInst_1_U2 ( .A(FSMReg[1]), .ZN(FSMMUX_MUXInst_1_n4) );
  NOR2_X1 FSMMUX_MUXInst_1_U1 ( .A1(rst), .A2(FSMMUX_MUXInst_1_n4), .ZN(
        FSMF[5]) );
  INV_X1 FSMMUX_MUXInst_2_U2 ( .A(FSMReg[2]), .ZN(FSMMUX_MUXInst_2_n4) );
  NOR2_X1 FSMMUX_MUXInst_2_U1 ( .A1(rst), .A2(FSMMUX_MUXInst_2_n4), .ZN(
        FSMF[6]) );
  OR2_X1 FSMMUX_MUXInst_3_U1 ( .A1(FSMReg[3]), .A2(rst), .ZN(FSM[3]) );
  INV_X1 FSMMUX_MUXInst_4_U2 ( .A(FSMReg[4]), .ZN(FSMMUX_MUXInst_4_n4) );
  NOR2_X1 FSMMUX_MUXInst_4_U1 ( .A1(rst), .A2(FSMMUX_MUXInst_4_n4), .ZN(FSM[4]) );
  INV_X1 FSMMUX_MUXInst_5_U2 ( .A(FSMReg[5]), .ZN(FSMMUX_MUXInst_5_n4) );
  NOR2_X1 FSMMUX_MUXInst_5_U1 ( .A1(rst), .A2(FSMMUX_MUXInst_5_n4), .ZN(FSM[5]) );
  INV_X1 FSMMUX_MUXInst_6_U2 ( .A(FSMReg[6]), .ZN(FSMMUX_MUXInst_6_n4) );
  NOR2_X1 FSMMUX_MUXInst_6_U1 ( .A1(rst), .A2(FSMMUX_MUXInst_6_n4), .ZN(FSM[6]) );
  XNOR2_X1 F_FSM_Inst_LFInst_0_LFInst_0_U2 ( .A(
        F_FSM_Inst_LFInst_0_LFInst_0_n3), .B(FSMF[6]), .ZN(FSMF[0]) );
  XNOR2_X1 F_FSM_Inst_LFInst_0_LFInst_0_U1 ( .A(FSMF[3]), .B(FSMF[5]), .ZN(
        F_FSM_Inst_LFInst_0_LFInst_0_n3) );
  XOR2_X1 F_FSM_Inst_LFInst_0_LFInst_1_U1 ( .A(FSMF[5]), .B(FSMF[3]), .Z(
        FSMF[1]) );
  XOR2_X1 F_FSM_Inst_LFInst_0_LFInst_2_U1 ( .A(FSMF[3]), .B(FSMF[6]), .Z(
        FSMF[2]) );
  XOR2_X1 F_FSM_Inst_LFInst_0_LFInst_4_U1 ( .A(FSMF[5]), .B(FSMF[6]), .Z(
        FSMF[4]) );
  XNOR2_X1 F_FSM_Inst_LFInst_1_LFInst_0_U2 ( .A(
        F_FSM_Inst_LFInst_1_LFInst_0_n3), .B(FSM[5]), .ZN(FSMF[7]) );
  XNOR2_X1 F_FSM_Inst_LFInst_1_LFInst_0_U1 ( .A(FSM[3]), .B(FSM[4]), .ZN(
        F_FSM_Inst_LFInst_1_LFInst_0_n3) );
  XNOR2_X1 F_FSM_Inst_LFInst_1_LFInst_1_U2 ( .A(
        F_FSM_Inst_LFInst_1_LFInst_1_n3), .B(FSM[6]), .ZN(FSMF[8]) );
  XNOR2_X1 F_FSM_Inst_LFInst_1_LFInst_1_U1 ( .A(FSM[3]), .B(FSM[4]), .ZN(
        F_FSM_Inst_LFInst_1_LFInst_1_n3) );
  XOR2_X1 F_FSM_Inst_LFInst_1_LFInst_2_U1 ( .A(FSM[3]), .B(FSM[5]), .Z(FSMF[9]) );
  XOR2_X1 F_FSM_Inst_LFInst_1_LFInst_3_U1 ( .A(FSM[3]), .B(FSM[6]), .Z(
        FSMF[10]) );
  XOR2_X1 F_FSM_Inst_LFInst_1_LFInst_4_U1 ( .A(FSM[4]), .B(FSM[5]), .Z(
        FSMF[11]) );
  XOR2_X1 F_FSM_Inst_LFInst_1_LFInst_5_U1 ( .A(FSM[4]), .B(FSM[6]), .Z(
        FSMF[12]) );
  XOR2_X1 F_FSM_Inst_LFInst_1_LFInst_6_U1 ( .A(FSM[5]), .B(FSM[6]), .Z(
        FSMF[13]) );
  XOR2_X1 FSMErrorVecGen_XORInst_0_0_U1 ( .A(FSMF[0]), .B(Red_RoundConstant[0]), .Z(FSMErrorVec[0]) );
  XOR2_X1 FSMErrorVecGen_XORInst_0_1_U1 ( .A(FSMF[1]), .B(Red_RoundConstant[1]), .Z(FSMErrorVec[1]) );
  XOR2_X1 FSMErrorVecGen_XORInst_0_2_U1 ( .A(FSMF[2]), .B(Red_RoundConstant[2]), .Z(FSMErrorVec[2]) );
  XOR2_X1 FSMErrorVecGen_XORInst_0_3_U1 ( .A(FSMF[3]), .B(Red_RoundConstant[3]), .Z(FSMErrorVec[3]) );
  XOR2_X1 FSMErrorVecGen_XORInst_0_4_U1 ( .A(FSMF[4]), .B(Red_RoundConstant[4]), .Z(FSMErrorVec[4]) );
  XOR2_X1 FSMErrorVecGen_XORInst_0_5_U1 ( .A(FSMF[5]), .B(Red_RoundConstant[5]), .Z(FSMErrorVec[5]) );
  XOR2_X1 FSMErrorVecGen_XORInst_0_6_U1 ( .A(FSMF[6]), .B(Red_RoundConstant[6]), .Z(FSMErrorVec[6]) );
  XOR2_X1 FSMErrorVecGen_XORInst_1_0_U1 ( .A(FSMF[7]), .B(Red_RoundConstant[7]), .Z(FSMErrorVec[7]) );
  XOR2_X1 FSMErrorVecGen_XORInst_1_1_U1 ( .A(FSMF[8]), .B(Red_RoundConstant[8]), .Z(FSMErrorVec[8]) );
  XOR2_X2 FSMErrorVecGen_XORInst_1_2_U1 ( .A(FSMF[9]), .B(Red_RoundConstant[9]), .Z(FSMErrorVec[9]) );
  XOR2_X1 FSMErrorVecGen_XORInst_1_3_U1 ( .A(FSMF[10]), .B(
        Red_RoundConstant[10]), .Z(FSMErrorVec[10]) );
  XOR2_X1 FSMErrorVecGen_XORInst_1_4_U1 ( .A(FSMF[11]), .B(
        Red_RoundConstant[11]), .Z(FSMErrorVec[11]) );
  XOR2_X2 FSMErrorVecGen_XORInst_1_5_U1 ( .A(FSMF[12]), .B(
        Red_RoundConstant[12]), .Z(FSMErrorVec[12]) );
  XOR2_X1 FSMErrorVecGen_XORInst_1_6_U1 ( .A(FSMF[13]), .B(
        Red_RoundConstant[13]), .Z(FSMErrorVec[13]) );
  NOR4_X1 F_SD1_StateUpdate_Done_Inst_U4 ( .A1(RoundConstant[4]), .A2(
        RoundConstant[5]), .A3(RoundConstant[7]), .A4(RoundConstant[0]), .ZN(
        F_SD1_StateUpdate_Done_Inst_n5) );
  AND4_X2 F_SD1_StateUpdate_Done_Inst_U2 ( .A1(RoundConstant[6]), .A2(
        RoundConstant[1]), .A3(RoundConstant[2]), .A4(
        F_SD1_StateUpdate_Done_Inst_n5), .ZN(done) );
  XNOR2_X1 F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_0_U12 ( .A(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_0_n12), .B(
        FSMF[5]), .ZN(RoundConstant[1]) );
  AOI22_X1 F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_0_U11 ( .A1(
        FSMErrorVec[5]), .A2(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_0_n6), .B1(
        FSMErrorVec[4]), .B2(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_0_n11), .ZN(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_0_n12) );
  OAI21_X1 F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_0_U10 ( .B1(
        FSMErrorVec[2]), .B2(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_0_n8), .A(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_0_n10), .ZN(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_0_n11) );
  NAND3_X1 F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_0_U9 ( .A1(
        FSMErrorVec[2]), .A2(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_0_n9), .A3(
        FSMErrorVec[5]), .ZN(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_0_n10) );
  NOR2_X1 F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_0_U8 ( .A1(
        FSMErrorVec[1]), .A2(FSMErrorVec[6]), .ZN(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_0_n9) );
  NOR3_X1 F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_0_U6 ( .A1(
        FSMErrorVec[3]), .A2(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_0_n4), .A3(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_0_n5), .ZN(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_0_n6) );
  INV_X1 F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_0_U5 ( .A(
        FSMErrorVec[1]), .ZN(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_0_n5) );
  NOR3_X1 F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_0_U4 ( .A1(
        FSMErrorVec[4]), .A2(FSMErrorVec[0]), .A3(FSMErrorVec[2]), .ZN(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_0_n4) );
  OAI33_X1 F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_0_U3 ( .A1(
        1'b0), .A2(FSMErrorVec[0]), .A3(1'b0), .B1(FSMErrorVec[5]), .B2(
        FSMErrorVec[1]), .B3(FSMErrorVec[3]), .ZN(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_0_n8) );
  XNOR2_X1 F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_1_U16 ( .A(
        FSMF[6]), .B(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_1_n13), .ZN(
        RoundConstant[2]) );
  AOI22_X1 F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_1_U15 ( .A1(
        FSMErrorVec[2]), .A2(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_1_n12), .B1(
        FSMErrorVec[6]), .B2(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_1_n11), .ZN(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_1_n13) );
  OAI22_X1 F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_1_U14 ( .A1(
        FSMErrorVec[5]), .A2(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_1_n10), .B1(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_1_n9), .B2(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_1_n8), .ZN(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_1_n11) );
  INV_X1 F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_1_U13 ( .A(
        FSMErrorVec[2]), .ZN(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_1_n8) );
  AOI21_X1 F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_1_U12 ( .B1(
        FSMErrorVec[1]), .B2(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_1_n7), .A(
        FSMErrorVec[4]), .ZN(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_1_n9) );
  AOI22_X1 F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_1_U11 ( .A1(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_1_n6), .A2(
        FSMErrorVec[2]), .B1(FSMErrorVec[4]), .B2(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_1_n5), .ZN(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_1_n10) );
  INV_X1 F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_1_U10 ( .A(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_1_n4), .ZN(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_1_n5) );
  AOI21_X1 F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_1_U9 ( .B1(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_1_n7), .B2(
        FSMErrorVec[0]), .A(FSMErrorVec[1]), .ZN(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_1_n4) );
  INV_X1 F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_1_U8 ( .A(
        FSMErrorVec[3]), .ZN(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_1_n7) );
  INV_X1 F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_1_U7 ( .A(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_1_n3), .ZN(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_1_n12) );
  OAI21_X1 F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_1_U6 ( .B1(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_1_n6), .B2(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_1_n2), .A(
        FSMErrorVec[4]), .ZN(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_1_n3) );
  AND3_X1 F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_1_U5 ( .A1(
        FSMErrorVec[1]), .A2(FSMErrorVec[5]), .A3(FSMErrorVec[3]), .ZN(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_1_n2) );
  NOR2_X1 F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_1_U4 ( .A1(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_1_n1), .A2(
        FSMErrorVec[1]), .ZN(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_1_n6) );
  INV_X1 F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_1_U3 ( .A(
        FSMErrorVec[0]), .ZN(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_1_n1) );
  XNOR2_X1 F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_2_U19 ( .A(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_2_n15), .B(
        RoundConstant[0]), .ZN(FSMUpdate[2]) );
  XOR2_X1 F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_2_U18 ( .A(
        FSMF[5]), .B(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_2_n14), .Z(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_2_n15) );
  AOI22_X1 F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_2_U17 ( .A1(
        FSMErrorVec[5]), .A2(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_2_n13), .B1(
        FSMErrorVec[4]), .B2(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_2_n12), .ZN(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_2_n14) );
  OAI22_X1 F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_2_U16 ( .A1(
        FSMErrorVec[2]), .A2(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_2_n11), .B1(
        FSMErrorVec[6]), .B2(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_2_n10), .ZN(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_2_n12) );
  NOR2_X1 F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_2_U15 ( .A1(
        FSMErrorVec[3]), .A2(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_2_n9), .ZN(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_2_n13) );
  XNOR2_X1 F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_2_U14 ( .A(
        FSMF[3]), .B(F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_2_n8), .ZN(RoundConstant[0]) );
  AOI22_X1 F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_2_U13 ( .A1(
        FSMErrorVec[3]), .A2(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_2_n7), .B1(
        FSMErrorVec[2]), .B2(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_2_n6), .ZN(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_2_n8) );
  NOR2_X1 F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_2_U12 ( .A1(
        FSMErrorVec[4]), .A2(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_2_n11), .ZN(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_2_n6) );
  OAI21_X1 F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_2_U11 ( .B1(
        FSMErrorVec[5]), .B2(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_2_n9), .A(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_2_n10), .ZN(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_2_n7) );
  NAND3_X1 F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_2_U10 ( .A1(
        FSMErrorVec[5]), .A2(FSMErrorVec[2]), .A3(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_2_n5), .ZN(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_2_n10) );
  INV_X1 F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_2_U9 ( .A(
        FSMErrorVec[1]), .ZN(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_2_n5) );
  INV_X1 F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_2_U7 ( .A(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_2_n5), .ZN(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_2_n3) );
  OAI21_X1 F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_2_U6 ( .B1(
        FSMErrorVec[3]), .B2(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_2_n2), .A(
        FSMErrorVec[0]), .ZN(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_2_n11) );
  NAND2_X1 F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_2_U5 ( .A1(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_2_n1), .A2(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_2_n5), .ZN(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_2_n2) );
  INV_X1 F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_2_U4 ( .A(
        FSMErrorVec[5]), .ZN(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_2_n1) );
  OAI33_X1 F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_2_U3 ( .A1(
        1'b0), .A2(F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_2_n3), 
        .A3(1'b0), .B1(FSMErrorVec[0]), .B2(FSMErrorVec[2]), .B3(
        FSMErrorVec[4]), .ZN(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_2_n9) );
  XNOR2_X1 F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_inst_3_U14 ( 
        .A(FSM[4]), .B(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_inst_3_n14), .ZN(
        RoundConstant[5]) );
  AOI22_X1 F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_inst_3_U13 ( 
        .A1(FSMErrorVec[12]), .A2(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_inst_3_n13), .B1(
        FSMErrorVec[11]), .B2(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_inst_3_n12), .ZN(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_inst_3_n14) );
  OAI21_X1 F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_inst_3_U12 ( 
        .B1(FSMErrorVec[9]), .B2(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_inst_3_n11), .A(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_inst_3_n10), .ZN(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_inst_3_n12) );
  NAND3_X1 F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_inst_3_U11 ( 
        .A1(FSMErrorVec[9]), .A2(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_inst_3_n9), .A3(
        FSMErrorVec[12]), .ZN(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_inst_3_n10) );
  NOR2_X1 F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_inst_3_U10 ( 
        .A1(FSMErrorVec[8]), .A2(FSMErrorVec[13]), .ZN(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_inst_3_n9) );
  NOR3_X1 F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_inst_3_U9 ( 
        .A1(FSMErrorVec[10]), .A2(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_inst_3_n8), .A3(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_inst_3_n5), .ZN(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_inst_3_n13) );
  NOR3_X1 F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_inst_3_U8 ( 
        .A1(FSMErrorVec[7]), .A2(FSMErrorVec[9]), .A3(FSMErrorVec[11]), .ZN(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_inst_3_n8) );
  INV_X1 F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_inst_3_U7 ( .A(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_inst_3_n7), .ZN(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_inst_3_n11) );
  INV_X1 F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_inst_3_U6 ( .A(
        FSMErrorVec[7]), .ZN(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_inst_3_n6) );
  INV_X1 F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_inst_3_U5 ( .A(
        FSMErrorVec[8]), .ZN(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_inst_3_n5) );
  NOR2_X1 F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_inst_3_U4 ( 
        .A1(FSMErrorVec[10]), .A2(FSMErrorVec[12]), .ZN(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_inst_3_n4) );
  AOI21_X1 F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_inst_3_U3 ( 
        .B1(F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_inst_3_n4), 
        .B2(F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_inst_3_n5), 
        .A(F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_inst_3_n6), 
        .ZN(F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_inst_3_n7) );
  INV_X1 F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_inst_4_U15 ( .A(
        FSMErrorVec[10]), .ZN(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_inst_4_n1) );
  XNOR2_X1 F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_inst_4_U14 ( 
        .A(F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_inst_4_n12), 
        .B(FSM[5]), .ZN(RoundConstant[6]) );
  AOI22_X1 F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_inst_4_U13 ( 
        .A1(FSMErrorVec[13]), .A2(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_inst_4_n4), .B1(
        FSMErrorVec[9]), .B2(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_inst_4_n11), .ZN(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_inst_4_n12) );
  OAI21_X1 F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_inst_4_U12 ( 
        .B1(F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_inst_4_n6), 
        .B2(F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_inst_4_n3), 
        .A(F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_inst_4_n10), 
        .ZN(F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_inst_4_n11)
         );
  OAI21_X1 F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_inst_4_U11 ( 
        .B1(FSMErrorVec[11]), .B2(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_inst_4_n9), .A(
        FSMErrorVec[13]), .ZN(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_inst_4_n10) );
  INV_X1 F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_inst_4_U9 ( .A(
        FSMErrorVec[7]), .ZN(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_inst_4_n7) );
  OAI222_X1 F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_inst_4_U8 ( 
        .A1(F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_inst_4_n5), 
        .A2(FSMErrorVec[10]), .B1(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_inst_4_n5), .B2(
        FSMErrorVec[12]), .C1(FSMErrorVec[7]), .C2(FSMErrorVec[8]), .ZN(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_inst_4_n6) );
  INV_X1 F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_inst_4_U7 ( .A(
        FSMErrorVec[8]), .ZN(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_inst_4_n5) );
  NOR3_X1 F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_inst_4_U6 ( 
        .A1(FSMErrorVec[12]), .A2(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_inst_4_n2), .A3(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_inst_4_n3), .ZN(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_inst_4_n4) );
  INV_X1 F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_inst_4_U5 ( .A(
        FSMErrorVec[11]), .ZN(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_inst_4_n3) );
  AOI21_X1 F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_inst_4_U4 ( 
        .B1(FSMErrorVec[7]), .B2(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_inst_4_n1), .A(
        FSMErrorVec[8]), .ZN(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_inst_4_n2) );
  OAI33_X1 F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_inst_4_U3 ( 
        .A1(1'b0), .A2(FSMErrorVec[10]), .A3(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_inst_4_n5), .B1(
        FSMErrorVec[8]), .B2(FSMErrorVec[12]), .B3(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_inst_4_n7), .ZN(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_inst_4_n9) );
  XOR2_X1 F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_inst_5_U15 ( 
        .A(FSM[6]), .B(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_inst_5_n12), .Z(
        RoundConstant[7]) );
  OAI21_X1 F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_inst_5_U14 ( 
        .B1(F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_inst_5_n11), 
        .B2(F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_inst_5_n10), 
        .A(F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_inst_5_n9), 
        .ZN(F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_inst_5_n12)
         );
  OAI211_X1 F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_inst_5_U13 ( 
        .C1(FSMErrorVec[12]), .C2(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_inst_5_n8), .A(
        FSMErrorVec[10]), .B(FSMErrorVec[13]), .ZN(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_inst_5_n9) );
  AOI221_X1 F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_inst_5_U12 ( 
        .B1(FSMErrorVec[8]), .B2(FSMErrorVec[11]), .C1(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_inst_5_n7), .C2(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_inst_5_n6), .A(
        FSMErrorVec[9]), .ZN(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_inst_5_n8) );
  AOI22_X1 F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_inst_5_U11 ( 
        .A1(F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_inst_5_n5), 
        .A2(F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_inst_5_n4), 
        .B1(FSMErrorVec[8]), .B2(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_inst_5_n3), .ZN(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_inst_5_n10) );
  AOI221_X1 F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_inst_5_U10 ( 
        .B1(F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_inst_5_n6), 
        .B2(FSMErrorVec[7]), .C1(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_inst_5_n2), .C2(
        FSMErrorVec[7]), .A(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_inst_5_n1), .ZN(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_inst_5_n3) );
  INV_X1 F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_inst_5_U9 ( .A(
        FSMErrorVec[10]), .ZN(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_inst_5_n1) );
  INV_X1 F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_inst_5_U8 ( .A(
        FSMErrorVec[9]), .ZN(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_inst_5_n2) );
  XNOR2_X1 F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_inst_5_U7 ( 
        .A(FSMErrorVec[9]), .B(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_inst_5_n7), .ZN(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_inst_5_n4) );
  INV_X1 F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_inst_5_U6 ( .A(
        FSMErrorVec[8]), .ZN(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_inst_5_n7) );
  AND2_X1 F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_inst_5_U5 ( 
        .A1(F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_inst_5_n6), 
        .A2(FSMErrorVec[13]), .ZN(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_inst_5_n5) );
  INV_X1 F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_inst_5_U4 ( .A(
        FSMErrorVec[11]), .ZN(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_inst_5_n6) );
  INV_X1 F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_inst_5_U3 ( .A(
        FSMErrorVec[12]), .ZN(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_inst_5_n11) );
  XNOR2_X1 F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_6_U21 ( .A(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_6_n17), .B(
        RoundConstant[4]), .ZN(FSMUpdate[6]) );
  XOR2_X1 F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_6_U20 ( .A(
        FSM[4]), .B(F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_6_n16), .Z(F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_6_n17) );
  AOI22_X1 F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_6_U19 ( .A1(
        FSMErrorVec[12]), .A2(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_6_n15), .B1(
        FSMErrorVec[11]), .B2(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_6_n14), .ZN(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_6_n16) );
  OAI22_X1 F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_6_U18 ( .A1(
        FSMErrorVec[9]), .A2(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_6_n13), .B1(
        FSMErrorVec[13]), .B2(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_6_n12), .ZN(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_6_n14) );
  NOR2_X1 F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_6_U17 ( .A1(
        FSMErrorVec[10]), .A2(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_6_n11), .ZN(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_6_n15) );
  XNOR2_X1 F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_6_U16 ( .A(
        FSM[3]), .B(F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_6_n10), .ZN(RoundConstant[4]) );
  AOI22_X1 F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_6_U15 ( .A1(
        FSMErrorVec[10]), .A2(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_6_n9), .B1(
        FSMErrorVec[9]), .B2(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_6_n8), .ZN(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_6_n10) );
  NOR2_X1 F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_6_U14 ( .A1(
        FSMErrorVec[11]), .A2(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_6_n13), .ZN(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_6_n8) );
  OAI21_X1 F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_6_U13 ( .B1(
        FSMErrorVec[12]), .B2(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_6_n11), .A(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_6_n12), .ZN(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_6_n9) );
  NAND3_X1 F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_6_U12 ( .A1(
        FSMErrorVec[12]), .A2(FSMErrorVec[9]), .A3(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_6_n2), .ZN(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_6_n12) );
  INV_X1 F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_6_U11 ( .A(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_6_n7), .ZN(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_6_n11) );
  INV_X1 F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_6_U10 ( .A(
        FSMErrorVec[9]), .ZN(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_6_n6) );
  INV_X1 F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_6_U9 ( .A(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_6_n4), .ZN(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_6_n13) );
  INV_X1 F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_6_U8 ( .A(
        FSMErrorVec[7]), .ZN(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_6_n3) );
  INV_X1 F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_6_U7 ( .A(
        FSMErrorVec[8]), .ZN(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_6_n2) );
  NOR2_X1 F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_6_U6 ( .A1(
        FSMErrorVec[11]), .A2(FSMErrorVec[7]), .ZN(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_6_n5) );
  AOI21_X1 F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_6_U5 ( .B1(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_6_n5), .B2(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_6_n6), .A(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_6_n2), .ZN(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_6_n7) );
  NOR2_X1 F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_6_U4 ( .A1(
        FSMErrorVec[12]), .A2(FSMErrorVec[10]), .ZN(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_6_n1) );
  AOI21_X1 F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_6_U3 ( .B1(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_6_n1), .B2(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_6_n2), .A(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_6_n3), .ZN(
        F_SD1_StateUpdate_Done_Inst_SD1_StateUpdate_Done_bit_6_n4) );
  DFF_X1 FSMRegInst_s_current_state_reg_0_ ( .D(RoundConstant[1]), .CK(clk), 
        .Q(FSMReg[0]), .QN() );
  DFF_X1 FSMRegInst_s_current_state_reg_1_ ( .D(RoundConstant[2]), .CK(clk), 
        .Q(FSMReg[1]), .QN() );
  DFF_X1 FSMRegInst_s_current_state_reg_2_ ( .D(FSMUpdate[2]), .CK(clk), .Q(
        FSMReg[2]), .QN() );
  DFF_X1 FSMRegInst_s_current_state_reg_3_ ( .D(RoundConstant[5]), .CK(clk), 
        .Q(FSMReg[3]), .QN() );
  DFF_X1 FSMRegInst_s_current_state_reg_4_ ( .D(RoundConstant[6]), .CK(clk), 
        .Q(FSMReg[4]), .QN() );
  DFF_X1 FSMRegInst_s_current_state_reg_5_ ( .D(RoundConstant[7]), .CK(clk), 
        .Q(FSMReg[5]), .QN() );
  DFF_X1 FSMRegInst_s_current_state_reg_6_ ( .D(FSMUpdate[6]), .CK(clk), .Q(
        FSMReg[6]), .QN() );
  NOR2_X1 selectsMUX_MUXInst_0_U1 ( .A1(selectsReg_0_), .A2(rst), .ZN(
        KeyMux_sel_input[4]) );
  INV_X1 F_SD1_SelectsUpdate_Bit0_Inst_U12 ( .A(
        F_SD1_SelectsUpdate_Bit0_Inst_n11), .ZN(selectsNext_0_) );
  OAI21_X1 F_SD1_SelectsUpdate_Bit0_Inst_U11 ( .B1(
        F_SD1_SelectsUpdate_Bit0_Inst_n10), .B2(
        F_SD1_SelectsUpdate_Bit0_Inst_n9), .A(F_SD1_SelectsUpdate_Bit0_Inst_n8), .ZN(F_SD1_SelectsUpdate_Bit0_Inst_n11) );
  NAND3_X1 F_SD1_SelectsUpdate_Bit0_Inst_U10 ( .A1(
        F_SD1_SelectsUpdate_Bit0_Inst_n7), .A2(n7), .A3(n4), .ZN(
        F_SD1_SelectsUpdate_Bit0_Inst_n8) );
  NOR3_X1 F_SD1_SelectsUpdate_Bit0_Inst_U9 ( .A1(
        F_SD1_SelectsUpdate_Bit0_Inst_n7), .A2(n7), .A3(n4), .ZN(
        F_SD1_SelectsUpdate_Bit0_Inst_n9) );
  XNOR2_X1 F_SD1_SelectsUpdate_Bit0_Inst_U8 ( .A(n3), .B(
        F_SD1_SelectsUpdate_Bit0_Inst_n6), .ZN(
        F_SD1_SelectsUpdate_Bit0_Inst_n7) );
  AOI21_X1 F_SD1_SelectsUpdate_Bit0_Inst_U7 ( .B1(n6), .B2(n5), .A(
        F_SD1_SelectsUpdate_Bit0_Inst_n5), .ZN(
        F_SD1_SelectsUpdate_Bit0_Inst_n10) );
  NOR2_X1 F_SD1_SelectsUpdate_Bit0_Inst_U6 ( .A1(
        F_SD1_SelectsUpdate_Bit0_Inst_n6), .A2(
        F_SD1_SelectsUpdate_Bit0_Inst_n3), .ZN(
        F_SD1_SelectsUpdate_Bit0_Inst_n5) );
  OAI21_X1 F_SD1_SelectsUpdate_Bit0_Inst_U5 ( .B1(n5), .B2(n6), .A(
        F_SD1_SelectsUpdate_Bit0_Inst_n4), .ZN(
        F_SD1_SelectsUpdate_Bit0_Inst_n6) );
  NAND2_X1 F_SD1_SelectsUpdate_Bit0_Inst_U4 ( .A1(n5), .A2(n6), .ZN(
        F_SD1_SelectsUpdate_Bit0_Inst_n4) );
  INV_X1 F_SD1_SelectsUpdate_Bit0_Inst_U3 ( .A(n3), .ZN(
        F_SD1_SelectsUpdate_Bit0_Inst_n3) );
  DFF_X1 selectsRegInst_s_current_state_reg_0_ ( .D(selectsNext_0_), .CK(clk), 
        .Q(), .QN(selectsReg_0_) );
  OR2_X1 Red_FSMMUX_MUXInst_0_U1 ( .A1(Red_FSMReg[0]), .A2(rst), .ZN(
        Red_RoundConstant[0]) );
  OR2_X1 Red_FSMMUX_MUXInst_1_U1 ( .A1(Red_FSMReg[1]), .A2(rst), .ZN(
        Red_RoundConstant[1]) );
  OR2_X1 Red_FSMMUX_MUXInst_2_U1 ( .A1(Red_FSMReg[2]), .A2(rst), .ZN(
        Red_RoundConstant[2]) );
  OR2_X1 Red_FSMMUX_MUXInst_3_U1 ( .A1(Red_FSMReg[3]), .A2(rst), .ZN(
        Red_RoundConstant[3]) );
  INV_X1 Red_FSMMUX_MUXInst_4_U2 ( .A(Red_FSMReg[4]), .ZN(
        Red_FSMMUX_MUXInst_4_n4) );
  NOR2_X2 Red_FSMMUX_MUXInst_4_U1 ( .A1(rst), .A2(Red_FSMMUX_MUXInst_4_n4), 
        .ZN(Red_RoundConstant[4]) );
  INV_X1 Red_FSMMUX_MUXInst_5_U2 ( .A(Red_FSMReg[5]), .ZN(
        Red_FSMMUX_MUXInst_5_n4) );
  NOR2_X2 Red_FSMMUX_MUXInst_5_U1 ( .A1(rst), .A2(Red_FSMMUX_MUXInst_5_n4), 
        .ZN(Red_RoundConstant[5]) );
  INV_X1 Red_FSMMUX_MUXInst_6_U2 ( .A(Red_FSMReg[6]), .ZN(
        Red_FSMMUX_MUXInst_6_n4) );
  NOR2_X2 Red_FSMMUX_MUXInst_6_U1 ( .A1(rst), .A2(Red_FSMMUX_MUXInst_6_n4), 
        .ZN(Red_RoundConstant[6]) );
  OR2_X1 Red_FSMMUX_MUXInst_7_U1 ( .A1(Red_FSMReg[7]), .A2(rst), .ZN(
        Red_RoundConstant[7]) );
  OR2_X2 Red_FSMMUX_MUXInst_8_U1 ( .A1(Red_FSMReg[8]), .A2(rst), .ZN(
        Red_RoundConstant[8]) );
  OR2_X1 Red_FSMMUX_MUXInst_9_U1 ( .A1(Red_FSMReg[9]), .A2(rst), .ZN(
        Red_RoundConstant[9]) );
  OR2_X1 Red_FSMMUX_MUXInst_10_U1 ( .A1(Red_FSMReg[10]), .A2(rst), .ZN(
        Red_RoundConstant[10]) );
  INV_X1 Red_FSMMUX_MUXInst_11_U2 ( .A(Red_FSMReg[11]), .ZN(
        Red_FSMMUX_MUXInst_11_n4) );
  NOR2_X2 Red_FSMMUX_MUXInst_11_U1 ( .A1(rst), .A2(Red_FSMMUX_MUXInst_11_n4), 
        .ZN(Red_RoundConstant[11]) );
  INV_X1 Red_FSMMUX_MUXInst_12_U2 ( .A(Red_FSMReg[12]), .ZN(
        Red_FSMMUX_MUXInst_12_n4) );
  NOR2_X4 Red_FSMMUX_MUXInst_12_U1 ( .A1(rst), .A2(Red_FSMMUX_MUXInst_12_n4), 
        .ZN(Red_RoundConstant[12]) );
  INV_X1 Red_FSMMUX_MUXInst_13_U2 ( .A(Red_FSMReg[13]), .ZN(
        Red_FSMMUX_MUXInst_13_n4) );
  NOR2_X2 Red_FSMMUX_MUXInst_13_U1 ( .A1(rst), .A2(Red_FSMMUX_MUXInst_13_n4), 
        .ZN(Red_RoundConstant[13]) );
  BUF_X2 F_SD2_RedStateUpdate_Done_Inst_U7 ( .A(FSM[4]), .Z(
        F_SD2_RedStateUpdate_Done_Inst_n7) );
  BUF_X2 F_SD2_RedStateUpdate_Done_Inst_U6 ( .A(FSMF[3]), .Z(
        F_SD2_RedStateUpdate_Done_Inst_n3) );
  BUF_X2 F_SD2_RedStateUpdate_Done_Inst_U5 ( .A(FSM[5]), .Z(
        F_SD2_RedStateUpdate_Done_Inst_n8) );
  BUF_X2 F_SD2_RedStateUpdate_Done_Inst_U4 ( .A(FSM[6]), .Z(
        F_SD2_RedStateUpdate_Done_Inst_n9) );
  BUF_X2 F_SD2_RedStateUpdate_Done_Inst_U3 ( .A(FSM[3]), .Z(
        F_SD2_RedStateUpdate_Done_Inst_n6) );
  BUF_X2 F_SD2_RedStateUpdate_Done_Inst_U2 ( .A(FSMF[6]), .Z(
        F_SD2_RedStateUpdate_Done_Inst_n5) );
  BUF_X2 F_SD2_RedStateUpdate_Done_Inst_U1 ( .A(FSMF[5]), .Z(
        F_SD2_RedStateUpdate_Done_Inst_n4) );
  OAI211_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_U139 ( 
        .C1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n329), .C2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n328), .A(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n326), 
        .B(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n325), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n327) );
  AOI221_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_U138 ( 
        .B1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n324), .B2(Red_RoundConstant[7]), .C1(Red_RoundConstant[8]), .C2(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n323), .A(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n322), 
        .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n325) );
  OAI22_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_U137 ( 
        .A1(Red_RoundConstant[7]), .A2(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n324), .B1(Red_RoundConstant[8]), .B2(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n323), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n322) );
  AOI21_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_U136 ( 
        .B1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n321), .B2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n320), .A(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n319), 
        .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n323) );
  OAI211_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_U135 ( 
        .C1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n318), .C2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n317), .A(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n316), 
        .B(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n315), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n319) );
  NAND3_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_U134 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n314), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n313), .A3(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n312), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n315) );
  OAI22_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_U133 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n311), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n310), .B1(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n309), .B2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n308), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n316) );
  AND3_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_U132 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n311), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n310), .A3(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n307), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n308) );
  NOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_U131 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n314), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n306), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n310) );
  OAI221_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_U130 ( 
        .B1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n305), .B2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n304), .C1(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n305), .C2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n303), .A(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n306), 
        .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n318) );
  NAND2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_U129 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n302), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n301), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n324) );
  OAI221_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_U128 ( 
        .B1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n300), .B2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n299), .C1(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n300), .C2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n298), .A(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n306), 
        .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n301) );
  OAI221_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_U127 ( 
        .B1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n297), .B2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n304), .C1(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n297), .C2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n296), .A(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n295), 
        .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n302) );
  OAI22_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_U126 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n320), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n294), .B1(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n293), .B2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n298), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n296) );
  NAND2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_U125 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n303), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n312), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n294) );
  AND2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_U124 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n313), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n305), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n297) );
  NOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_U123 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n312), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n298), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n305) );
  AOI21_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_U122 ( 
        .B1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n292), .B2(Red_RoundConstant[9]), .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n291), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n326) );
  OAI211_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_U121 ( 
        .C1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n292), .C2(Red_RoundConstant[9]), .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n290), .B(Red_FSMUpdate[0]), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n291) );
  AOI221_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_U120 ( 
        .B1(Red_RoundConstant[0]), .B2(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n289), .C1(Red_RoundConstant[12]), .C2(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n288), .A(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n287), 
        .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n290) );
  OAI22_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_U119 ( 
        .A1(Red_RoundConstant[0]), .A2(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n289), .B1(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n288), .B2(Red_RoundConstant[12]), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n287) );
  AOI221_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_U118 ( 
        .B1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n286), .B2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n303), .C1(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n285), .C2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n303), .A(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n284), 
        .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n288) );
  AOI221_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_U117 ( 
        .B1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n304), .B2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n295), .C1(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n283), .C2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n282), .A(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n281), 
        .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n284) );
  OAI21_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_U116 ( 
        .B1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n306), .B2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n280), .A(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n279), 
        .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n285) );
  OAI21_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_U115 ( 
        .B1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n278), .B2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n298), .A(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n277), 
        .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n279) );
  INV_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_U114 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n276), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n277) );
  AOI21_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_U113 ( 
        .B1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n311), .B2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n320), .A(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n275), 
        .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n276) );
  AOI22_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_U112 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n311), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n293), .B1(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n274), .B2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n298), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n280) );
  NOR3_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_U111 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n304), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n314), .A3(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n298), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n286) );
  OAI211_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_U110 ( 
        .C1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n312), .C2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n258), .A(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n257), 
        .B(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n256), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n292) );
  OAI21_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_U109 ( 
        .B1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n300), .B2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n255), .A(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n275), 
        .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n256) );
  OAI22_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_U108 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n306), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n254), .B1(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n253), .B2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n252), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n255) );
  NAND2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_U107 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n303), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n293), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n252) );
  INV_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_U106 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n299), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n254) );
  NOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_U105 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n303), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n251), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n299) );
  NOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_U104 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n311), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n274), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n251) );
  INV_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_U103 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n250), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n300) );
  AOI21_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_U102 ( 
        .B1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n274), .B2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n311), .A(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n321), 
        .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n250) );
  NOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_U101 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n249), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n282), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n321) );
  NAND2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_U100 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n253), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n314), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n282) );
  INV_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_U99 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n293), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n314) );
  NOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_U98 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n304), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n253), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n311) );
  INV_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_U97 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n312), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n253) );
  INV_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_U96 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n317), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n274) );
  NAND2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_U95 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n320), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n293), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n317) );
  NAND4_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_U94 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n248), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n278), .A3(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n312), .A4(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n320), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n257) );
  NOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_U93 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n283), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n293), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n278) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_U92 ( 
        .A(Red_RoundConstant[13]), .B(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n247), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n293) );
  XOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_U91 ( 
        .A(F_SD2_RedStateUpdate_Done_Inst_n8), .B(
        F_SD2_RedStateUpdate_Done_Inst_n9), .Z(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n247) );
  INV_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_U90 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n304), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n283) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_U89 ( 
        .A(Red_RoundConstant[11]), .B(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n246), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n304) );
  NOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_U88 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n275), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n295), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n248) );
  NAND2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_U87 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n306), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n309), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n258) );
  INV_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_U86 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n281), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n309) );
  NAND2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_U85 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n298), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n313), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n281) );
  NOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_U84 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n320), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n303), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n313) );
  INV_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_U83 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n249), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n303) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_U82 ( 
        .A(Red_RoundConstant[12]), .B(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n245), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n249) );
  XOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_U81 ( 
        .A(F_SD2_RedStateUpdate_Done_Inst_n7), .B(
        F_SD2_RedStateUpdate_Done_Inst_n9), .Z(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n245) );
  INV_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_U80 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n307), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n320) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_U79 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n244), .B(Red_RoundConstant[8]), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n307) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_U78 ( 
        .A(F_SD2_RedStateUpdate_Done_Inst_n7), .B(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n243), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n244) );
  INV_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_U77 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n275), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n298) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_U76 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n242), .B(Red_RoundConstant[9]), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n275) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_U75 ( 
        .A(F_SD2_RedStateUpdate_Done_Inst_n8), .B(
        F_SD2_RedStateUpdate_Done_Inst_n6), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n242) );
  INV_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_U74 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n295), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n306) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_U73 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n241), .B(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n246), 
        .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n295) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_U72 ( 
        .A(F_SD2_RedStateUpdate_Done_Inst_n8), .B(
        F_SD2_RedStateUpdate_Done_Inst_n7), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n246) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_U71 ( 
        .A(Red_RoundConstant[7]), .B(F_SD2_RedStateUpdate_Done_Inst_n6), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n241) );
  XOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_U70 ( 
        .A(Red_RoundConstant[10]), .B(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n240), .Z(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n312)
         );
  INV_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_U69 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n243), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n240) );
  XOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_U68 ( 
        .A(F_SD2_RedStateUpdate_Done_Inst_n6), .B(
        F_SD2_RedStateUpdate_Done_Inst_n9), .Z(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n243) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_U67 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n239), .B(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n238), 
        .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n328) );
  AOI211_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_U66 ( 
        .C1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n260), .C2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n237), .A(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n236), 
        .B(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n235), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n238) );
  AOI21_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_U65 ( 
        .B1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n234), .B2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n233), .A(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n232), 
        .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n235) );
  OAI211_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_U64 ( 
        .C1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n234), .C2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n233), .A(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n260), 
        .B(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n259), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n232) );
  AOI21_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_U63 ( 
        .B1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n231), .B2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n230), .A(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n229), 
        .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n236) );
  NAND3_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_U62 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n263), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n265), .A3(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n264), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n230) );
  INV_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_U61 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n228), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n231) );
  INV_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_U60 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n227), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n237) );
  AOI21_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_U59 ( 
        .B1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n226), .B2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n225), .A(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n224), 
        .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n227) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_U58 ( 
        .A(Red_RoundConstant[1]), .B(Red_RoundConstant[5]), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n239) );
  OAI211_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_U57 ( 
        .C1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n223), .C2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n229), .A(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n222), 
        .B(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n221), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n329) );
  NAND3_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_U56 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n260), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n228), .A3(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n220), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n221) );
  AOI221_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_U55 ( 
        .B1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n224), .B2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n266), .C1(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n219), .C2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n266), .A(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n218), 
        .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n222) );
  OAI22_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_U54 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n266), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n273), .B1(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n217), .B2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n216), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n218) );
  NAND2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_U53 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n269), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n220), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n216) );
  INV_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_U52 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n272), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n269) );
  NAND2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_U51 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n259), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n263), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n217) );
  NOR3_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_U50 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n260), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n263), .A3(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n234), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n219) );
  NOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_U49 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n268), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n215), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n224) );
  INV_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_U48 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n226), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n223) );
  NAND2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_U47 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n268), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n215), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n226) );
  NAND2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_U46 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n272), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n234), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n215) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_U45 ( 
        .A(Red_RoundConstant[2]), .B(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n214), .ZN(Red_FSMUpdate[0]) );
  AOI211_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_U44 ( 
        .C1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n259), .C2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n213), .A(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n212), 
        .B(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n211), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n214) );
  NOR3_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_U43 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n229), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n261), .A3(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n272), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n211) );
  NAND2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_U42 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n266), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n271), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n229) );
  NOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_U41 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n259), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n260), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n271) );
  AOI21_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_U40 ( 
        .B1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n210), .B2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n209), .A(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n263), 
        .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n212) );
  NAND3_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_U39 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n265), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n228), .A3(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n225), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n209) );
  NOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_U38 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n266), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n259), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n225) );
  NOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_U37 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n264), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n272), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n228) );
  NAND3_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_U36 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n260), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n259), .A3(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n234), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n210) );
  OAI211_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_U35 ( 
        .C1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n267), .C2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n268), .A(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n273), 
        .B(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n208), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n213) );
  NAND3_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_U34 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n262), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n272), .A3(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n270), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n208) );
  NAND2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_U33 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n268), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n267), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n270) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_U32 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n207), .B(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n206), 
        .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n272) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_U31 ( 
        .A(F_SD2_RedStateUpdate_Done_Inst_n3), .B(Red_RoundConstant[0]), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n207) );
  NAND2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_U30 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n263), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n205), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n273) );
  NOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_U29 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n262), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n234), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n205) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_U28 ( 
        .A(Red_RoundConstant[5]), .B(F_SD2_RedStateUpdate_Done_Inst_n4), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n262) );
  INV_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_U27 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n261), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n263) );
  NAND2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_U26 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n261), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n264), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n268) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_U25 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n206), .B(Red_RoundConstant[4]), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n233) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_U24 ( 
        .A(F_SD2_RedStateUpdate_Done_Inst_n4), .B(
        F_SD2_RedStateUpdate_Done_Inst_n5), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n206) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_U23 ( 
        .A(F_SD2_RedStateUpdate_Done_Inst_n3), .B(Red_RoundConstant[3]), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n261) );
  INV_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_U22 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n220), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n267) );
  NOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_U21 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n266), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n265), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n220) );
  INV_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_U20 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n234), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n265) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_U19 ( 
        .A(F_SD2_RedStateUpdate_Done_Inst_n5), .B(Red_RoundConstant[6]), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n234) );
  XOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_U18 ( 
        .A(F_SD2_RedStateUpdate_Done_Inst_n3), .B(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n204), .Z(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n266)
         );
  XOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_U17 ( 
        .A(Red_RoundConstant[1]), .B(F_SD2_RedStateUpdate_Done_Inst_n4), .Z(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n204) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_U16 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n203), .B(F_SD2_RedStateUpdate_Done_Inst_n5), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n259) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_U15 ( 
        .A(F_SD2_RedStateUpdate_Done_Inst_n3), .B(Red_RoundConstant[2]), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n203) );
  INV_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_U14 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n233), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n264) );
  INV_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_U13 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n262), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n260) );
  AOI21_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_U12 ( 
        .B1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n329), .B2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n328), .A(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n327), 
        .ZN(Red_done[0]) );
  AOI211_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_U11 ( 
        .C1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n272), .C2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n199), .A(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n200), 
        .B(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n202), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n289) );
  AOI21_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_U10 ( 
        .B1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n273), .B2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n201), .A(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n272), 
        .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n202) );
  NAND2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_U9 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n271), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n270), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n201) );
  NOR3_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_U8 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n268), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n267), .A3(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n272), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n200) );
  OAI21_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_U7 ( 
        .B1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n264), .B2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n198), .A(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n197), 
        .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n199) );
  NAND2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_U6 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n265), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n259), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n198) );
  NAND2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_U5 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n266), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n196), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n197) );
  OAI33_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_U4 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n195), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n261), .A3(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n260), .B1(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n262), .B2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n263), .B3(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n264), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n196) );
  INV_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_U3 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n259), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_0_n195) );
  OAI21_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_U128 ( 
        .B1(Red_RoundConstant[8]), .B2(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n314), .A(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n313), 
        .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n315) );
  AOI211_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_U127 ( 
        .C1(Red_RoundConstant[8]), .C2(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n314), .A(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n312), 
        .B(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n311), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n313) );
  OAI221_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_U126 ( 
        .B1(Red_RoundConstant[12]), .B2(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n310), .C1(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n309), .C2(Red_RoundConstant[9]), .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n308), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n311) );
  AOI22_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_U125 ( 
        .A1(Red_RoundConstant[12]), .A2(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n310), .B1(Red_RoundConstant[9]), .B2(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n309), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n308) );
  OAI221_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_U124 ( 
        .B1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n307), .B2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n306), .C1(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n307), .C2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n305), .A(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n304), 
        .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n309) );
  OAI221_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_U123 ( 
        .B1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n303), .B2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n302), .C1(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n301), .C2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n300), .A(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n299), 
        .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n304) );
  NOR3_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_U122 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n298), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n297), .A3(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n296), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n302) );
  AOI22_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_U121 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n295), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n294), .B1(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n293), .B2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n301), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n305) );
  NOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_U120 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n292), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n291), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n293) );
  AOI221_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_U119 ( 
        .B1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n290), .B2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n289), .C1(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n288), .C2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n289), .A(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n287), 
        .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n310) );
  AOI21_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_U118 ( 
        .B1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n286), .B2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n294), .A(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n285), 
        .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n287) );
  OAI21_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_U117 ( 
        .B1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n284), .B2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n286), .A(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n300), 
        .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n285) );
  OAI21_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_U116 ( 
        .B1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n307), .B2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n296), .A(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n283), 
        .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n288) );
  AOI22_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_U115 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n282), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n281), .B1(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n307), .B2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n280), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n283) );
  INV_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_U114 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n279), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n280) );
  AOI22_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_U113 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n278), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n282), .B1(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n294), .B2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n277), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n279) );
  NOR3_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_U112 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n286), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n292), .A3(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n307), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n290) );
  AOI21_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_U111 ( 
        .B1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n276), .B2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n278), .A(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n275), 
        .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n314) );
  OAI211_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_U110 ( 
        .C1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n274), .C2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n294), .A(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n273), 
        .B(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n272), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n275) );
  NAND3_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_U109 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n271), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n292), .A3(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n301), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n272) );
  INV_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_U108 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n270), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n271) );
  OAI22_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_U107 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n282), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n281), .B1(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n300), .B2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n269), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n273) );
  AND3_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_U106 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n282), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n281), .A3(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n297), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n269) );
  NOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_U105 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n298), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n270), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n300) );
  NOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_U104 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n292), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n299), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n281) );
  INV_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_U103 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n294), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n299) );
  OAI221_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_U102 ( 
        .B1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n268), .B2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n303), .C1(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n268), .C2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n298), .A(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n277), 
        .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n274) );
  INV_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_U101 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n267), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n268) );
  OAI221_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_U100 ( 
        .B1(Red_RoundConstant[7]), .B2(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n266), .C1(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n265), .C2(Red_RoundConstant[2]), .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n264), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n316) );
  AOI22_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_U99 ( 
        .A1(Red_RoundConstant[7]), .A2(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n266), .B1(Red_RoundConstant[2]), .B2(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n265), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n264) );
  OAI211_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_U98 ( 
        .C1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n263), .C2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n262), .A(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n261), 
        .B(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n260), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n265) );
  NAND4_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_U97 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n259), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n258), .A3(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n257), .A4(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n256), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n260) );
  INV_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_U96 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n255), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n256) );
  OAI221_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_U95 ( 
        .B1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n254), .B2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n253), .C1(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n254), .C2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n252), .A(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n251), 
        .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n261) );
  AOI21_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_U94 ( 
        .B1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n250), .B2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n249), .A(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n248), 
        .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n254) );
  OAI21_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_U93 ( 
        .B1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n253), .B2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n252), .A(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n247), 
        .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n249) );
  INV_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_U92 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n246), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n263) );
  OAI21_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_U91 ( 
        .B1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n245), .B2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n294), .A(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n244), 
        .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n266) );
  OAI21_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_U90 ( 
        .B1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n243), .B2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n242), .A(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n294), 
        .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n244) );
  NOR3_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_U89 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n303), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n278), .A3(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n267), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n242) );
  NAND2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_U88 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n286), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n289), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n267) );
  AOI221_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_U87 ( 
        .B1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n301), .B2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n296), .C1(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n270), .C2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n296), .A(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n307), 
        .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n243) );
  NAND2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_U86 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n297), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n291), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n270) );
  INV_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_U85 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n289), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n291) );
  NAND2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_U84 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n286), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n292), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n296) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_U83 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n241), .B(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n240), 
        .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n294) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_U82 ( 
        .A(F_SD2_RedStateUpdate_Done_Inst_n7), .B(Red_RoundConstant[7]), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n241) );
  AOI21_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_U81 ( 
        .B1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n295), .B2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n307), .A(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n239), 
        .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n245) );
  INV_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_U80 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n306), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n239) );
  AOI21_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_U79 ( 
        .B1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n282), .B2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n277), .A(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n276), 
        .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n306) );
  AND2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_U78 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n289), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n284), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n276) );
  AND2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_U77 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n303), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n292), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n284) );
  INV_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_U76 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n298), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n307) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_U75 ( 
        .A(Red_RoundConstant[9]), .B(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n240), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n298) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_U74 ( 
        .A(F_SD2_RedStateUpdate_Done_Inst_n6), .B(
        F_SD2_RedStateUpdate_Done_Inst_n8), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n240) );
  NOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_U73 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n289), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n238), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n295) );
  NOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_U72 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n282), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n277), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n238) );
  NOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_U71 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n297), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n292), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n277) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_U70 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n237), .B(Red_RoundConstant[13]), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n292) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_U69 ( 
        .A(F_SD2_RedStateUpdate_Done_Inst_n9), .B(
        F_SD2_RedStateUpdate_Done_Inst_n8), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n237) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_U68 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n236), .B(F_SD2_RedStateUpdate_Done_Inst_n7), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n297) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_U67 ( 
        .A(Red_RoundConstant[8]), .B(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n235), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n236) );
  NOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_U66 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n303), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n286), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n282) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_U65 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n234), .B(Red_RoundConstant[11]), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n286) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_U64 ( 
        .A(F_SD2_RedStateUpdate_Done_Inst_n8), .B(
        F_SD2_RedStateUpdate_Done_Inst_n7), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n234) );
  INV_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_U63 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n301), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n303) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_U62 ( 
        .A(Red_RoundConstant[10]), .B(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n235), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n301) );
  XOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_U61 ( 
        .A(F_SD2_RedStateUpdate_Done_Inst_n6), .B(
        F_SD2_RedStateUpdate_Done_Inst_n9), .Z(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n235) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_U60 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n233), .B(Red_RoundConstant[12]), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n289) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_U59 ( 
        .A(F_SD2_RedStateUpdate_Done_Inst_n9), .B(
        F_SD2_RedStateUpdate_Done_Inst_n7), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n233) );
  XOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_U58 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n317), .B(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n312), 
        .Z(Red_FSMUpdate[1]) );
  NOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_U57 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n228), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n259), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n252) );
  NAND2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_U56 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n228), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n262), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n250) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_U55 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n225), .B(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n224), 
        .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n317) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_U54 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n223), .B(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n222), 
        .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n224) );
  AOI221_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_U53 ( 
        .B1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n229), .B2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n247), .C1(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n221), .C2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n220), .A(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n219), 
        .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n222) );
  OAI22_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_U52 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n218), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n217), .B1(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n216), .B2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n230), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n219) );
  NAND3_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_U51 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n259), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n215), .A3(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n247), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n230) );
  INV_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_U50 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n232), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n259) );
  AOI22_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_U49 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n228), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n258), .B1(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n251), .B2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n214), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n216) );
  OAI22_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_U48 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n248), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n213), .B1(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n228), .B2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n255), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n221) );
  NAND2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_U47 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n248), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n262), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n255) );
  INV_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_U46 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n220), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n247) );
  NOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_U45 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n212), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n211), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n229) );
  OAI21_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_U44 ( 
        .B1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n212), .B2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n210), .A(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n209), 
        .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n223) );
  OAI21_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_U43 ( 
        .B1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n226), .B2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n246), .A(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n208), 
        .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n209) );
  OAI21_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_U42 ( 
        .B1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n217), .B2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n211), .A(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n226), 
        .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n208) );
  NAND2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_U41 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n248), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n214), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n211) );
  OAI22_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_U40 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n212), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n227), .B1(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n232), .B2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n217), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n246) );
  NAND2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_U39 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n220), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n231), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n217) );
  NOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_U38 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n228), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n251), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n231) );
  INV_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_U37 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n212), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n228) );
  NAND2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_U36 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n248), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n251), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n227) );
  AOI22_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_U35 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n257), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n207), .B1(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n215), .B2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n206), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n210) );
  OAI21_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_U34 ( 
        .B1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n258), .B2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n205), .A(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n213), 
        .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n206) );
  NAND2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_U33 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n253), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n232), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n213) );
  INV_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_U32 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n251), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n205) );
  INV_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_U31 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n218), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n207) );
  AOI21_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_U30 ( 
        .B1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n215), .B2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n232), .A(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n253), 
        .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n218) );
  NOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_U29 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n258), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n214), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n253) );
  XOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_U28 ( 
        .A(F_SD2_RedStateUpdate_Done_Inst_n3), .B(Red_RoundConstant[3]), .Z(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n214) );
  INV_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_U27 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n226), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n258) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_U26 ( 
        .A(Red_RoundConstant[4]), .B(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n204), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n226) );
  XOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_U25 ( 
        .A(F_SD2_RedStateUpdate_Done_Inst_n4), .B(
        F_SD2_RedStateUpdate_Done_Inst_n5), .Z(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n204) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_U24 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n203), .B(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n202), 
        .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n232) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_U23 ( 
        .A(F_SD2_RedStateUpdate_Done_Inst_n5), .B(Red_RoundConstant[0]), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n203) );
  INV_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_U22 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n248), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n215) );
  XOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_U21 ( 
        .A(Red_RoundConstant[6]), .B(F_SD2_RedStateUpdate_Done_Inst_n5), .Z(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n248) );
  NOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_U20 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n251), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n220), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n257) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_U19 ( 
        .A(Red_RoundConstant[1]), .B(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n202), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n220) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_U18 ( 
        .A(F_SD2_RedStateUpdate_Done_Inst_n4), .B(
        F_SD2_RedStateUpdate_Done_Inst_n3), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n202) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_U17 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n201), .B(F_SD2_RedStateUpdate_Done_Inst_n3), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n251) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_U16 ( 
        .A(F_SD2_RedStateUpdate_Done_Inst_n5), .B(Red_RoundConstant[2]), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n201) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_U15 ( 
        .A(Red_RoundConstant[5]), .B(F_SD2_RedStateUpdate_Done_Inst_n4), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n212) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_U14 ( 
        .A(Red_RoundConstant[5]), .B(Red_RoundConstant[1]), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n225) );
  INV_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_U13 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n214), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n262) );
  INV_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_U12 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n297), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n278) );
  NOR3_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_U11 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n317), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n316), .A3(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n315), .ZN(Red_done[1]) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_U10 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n200), .B(Red_RoundConstant[0]), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n312) );
  AOI211_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_U9 ( 
        .C1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n232), .C2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n194), .A(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n196), 
        .B(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n199), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n200) );
  OAI22_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_U8 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n232), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n197), .B1(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n198), .B2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n230), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n199) );
  NOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_U7 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n253), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n231), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n198) );
  AOI21_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_U6 ( 
        .B1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n231), .B2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n253), .A(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n229), 
        .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n197) );
  NOR3_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_U5 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n247), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n262), .A3(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n195), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n196) );
  NAND2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_U4 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n252), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n251), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n195) );
  AOI221_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_U3 ( 
        .B1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n247), .B2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n227), .C1(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n250), .C2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n227), .A(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n226), 
        .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_1_n194) );
  INV_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_U42 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_n233), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_n232) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_U41 ( 
        .A(F_SD2_RedStateUpdate_Done_Inst_n5), .B(
        F_SD2_RedStateUpdate_Done_Inst_n4), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_n233) );
  INV_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_U40 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_n198), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_n213) );
  INV_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_U39 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_n221), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_n226) );
  INV_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_U38 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_n207), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_n217) );
  XOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_U37 ( 
        .A(Red_RoundConstant[1]), .B(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_n231), .Z(Red_FSMUpdate[2]) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_U36 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_n230), .B(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_n229), 
        .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_n231) );
  OAI21_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_U35 ( 
        .B1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_n195), .B2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_n220), .A(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_n210), 
        .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_n230) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_U34 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_n228), .B(Red_RoundConstant[5]), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_n229) );
  OAI21_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_U33 ( 
        .B1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_n208), .B2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_n214), .A(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_n227), 
        .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_n228) );
  INV_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_U32 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_n214), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_n216) );
  OAI21_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_U31 ( 
        .B1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_n226), .B2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_n217), .A(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_n225), 
        .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_n227) );
  NAND3_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_U30 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_n224), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_n223), .A3(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_n217), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_n225) );
  NAND2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_U29 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_n203), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_n202), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_n224) );
  NAND3_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_U28 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_n198), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_n201), .A3(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_n222), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_n223) );
  OAI22_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_U27 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_n196), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_n195), .B1(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_n200), .B2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_n205), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_n222) );
  OAI221_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_U26 ( 
        .B1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_n195), .B2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_n212), .C1(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_n211), .C2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_n212), .A(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_n200), 
        .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_n221) );
  INV_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_U25 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_n208), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_n209) );
  AOI21_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_U24 ( 
        .B1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_n212), .B2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_n200), .A(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_n219), 
        .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_n220) );
  OAI21_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_U23 ( 
        .B1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_n205), .B2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_n215), .A(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_n218), 
        .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_n219) );
  NAND3_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_U22 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_n205), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_n216), .A3(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_n217), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_n218) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_U21 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_n211), .B(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_n196), 
        .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_n215) );
  AOI22_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_U20 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_n213), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_n201), .B1(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_n200), .B2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_n196), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_n214) );
  NOR3_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_U19 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_n198), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_n211), .A3(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_n199), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_n212) );
  INV_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_U18 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_n201), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_n211) );
  OAI221_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_U17 ( 
        .B1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_n196), .B2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_n198), .C1(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_n199), .C2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_n202), .A(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_n209), 
        .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_n210) );
  NAND3_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_U16 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_n195), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_n205), .A3(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_n207), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_n208) );
  XOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_U15 ( 
        .A(F_SD2_RedStateUpdate_Done_Inst_n3), .B(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_n206), .Z(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_n207)
         );
  XOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_U14 ( 
        .A(F_SD2_RedStateUpdate_Done_Inst_n4), .B(Red_RoundConstant[1]), .Z(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_n206) );
  XOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_U13 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_n204), .B(Red_RoundConstant[2]), .Z(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_n205) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_U12 ( 
        .A(F_SD2_RedStateUpdate_Done_Inst_n5), .B(
        F_SD2_RedStateUpdate_Done_Inst_n3), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_n204) );
  INV_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_U11 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_n195), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_n203) );
  NOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_U10 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_n200), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_n201), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_n202) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_U9 ( 
        .A(F_SD2_RedStateUpdate_Done_Inst_n5), .B(Red_RoundConstant[6]), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_n201) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_U8 ( 
        .A(F_SD2_RedStateUpdate_Done_Inst_n3), .B(Red_RoundConstant[3]), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_n200) );
  INV_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_U7 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_n196), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_n199) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_U6 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_n197), .B(Red_RoundConstant[0]), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_n198) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_U5 ( 
        .A(F_SD2_RedStateUpdate_Done_Inst_n3), .B(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_n232), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_n197) );
  XOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_U4 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_n233), .B(Red_RoundConstant[4]), .Z(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_n196) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_U3 ( 
        .A(F_SD2_RedStateUpdate_Done_Inst_n4), .B(Red_RoundConstant[5]), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_2_n195) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_U38 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_n228), .B(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_n227), 
        .ZN(Red_FSMUpdate[3]) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_U37 ( 
        .A(Red_RoundConstant[0]), .B(Red_RoundConstant[2]), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_n227) );
  XOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_U36 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_n226), .B(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_n225), 
        .Z(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_n228) );
  OAI21_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_U35 ( 
        .B1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_n224), .B2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_n223), .A(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_n222), 
        .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_n225) );
  OAI21_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_U34 ( 
        .B1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_n221), .B2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_n220), .A(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_n224), 
        .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_n222) );
  OAI22_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_U33 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_n219), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_n218), .B1(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_n217), .B2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_n216), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_n221) );
  AOI21_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_U32 ( 
        .B1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_n215), .B2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_n214), .A(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_n213), 
        .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_n218) );
  AOI21_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_U31 ( 
        .B1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_n216), .B2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_n217), .A(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_n212), 
        .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_n213) );
  OR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_U30 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_n211), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_n215), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_n217) );
  OAI21_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_U29 ( 
        .B1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_n210), .B2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_n209), .A(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_n211), 
        .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_n223) );
  AND3_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_U28 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_n208), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_n207), .A3(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_n206), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_n209) );
  OAI21_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_U27 ( 
        .B1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_n205), .B2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_n211), .A(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_n204), 
        .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_n226) );
  OAI21_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_U26 ( 
        .B1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_n203), .B2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_n220), .A(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_n211), 
        .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_n204) );
  NOR3_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_U25 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_n208), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_n214), .A3(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_n202), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_n220) );
  AOI222_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_U24 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_n216), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_n201), .B1(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_n216), .B2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_n200), .C1(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_n201), .C2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_n200), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_n203) );
  OR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_U23 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_n215), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_n224), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_n200) );
  NAND2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_U22 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_n208), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_n199), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_n201) );
  NAND2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_U21 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_n207), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_n214), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_n216) );
  XOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_U20 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_n198), .B(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_n197), 
        .Z(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_n211) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_U19 ( 
        .A(Red_RoundConstant[0]), .B(F_SD2_RedStateUpdate_Done_Inst_n3), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_n198) );
  AOI221_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_U18 ( 
        .B1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_n210), .B2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_n224), .C1(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_n206), .C2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_n224), .A(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_n196), 
        .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_n205) );
  NOR4_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_U17 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_n219), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_n199), .A3(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_n207), .A4(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_n202), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_n196) );
  INV_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_U16 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_n215), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_n202) );
  NOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_U15 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_n199), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_n214), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_n206) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_U14 ( 
        .A(F_SD2_RedStateUpdate_Done_Inst_n5), .B(Red_RoundConstant[6]), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_n214) );
  INV_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_U13 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_n212), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_n199) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_U12 ( 
        .A(Red_RoundConstant[4]), .B(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_n197), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_n212) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_U11 ( 
        .A(F_SD2_RedStateUpdate_Done_Inst_n4), .B(
        F_SD2_RedStateUpdate_Done_Inst_n5), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_n197) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_U10 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_n195), .B(F_SD2_RedStateUpdate_Done_Inst_n5), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_n224) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_U9 ( 
        .A(Red_RoundConstant[2]), .B(F_SD2_RedStateUpdate_Done_Inst_n3), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_n195) );
  NOR3_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_U8 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_n215), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_n207), .A3(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_n208), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_n210) );
  INV_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_U7 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_n219), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_n208) );
  XOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_U6 ( 
        .A(F_SD2_RedStateUpdate_Done_Inst_n3), .B(Red_RoundConstant[3]), .Z(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_n219) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_U5 ( 
        .A(Red_RoundConstant[1]), .B(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_n194), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_n207) );
  XOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_U4 ( 
        .A(F_SD2_RedStateUpdate_Done_Inst_n3), .B(
        F_SD2_RedStateUpdate_Done_Inst_n4), .Z(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_n194) );
  XOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_U3 ( 
        .A(F_SD2_RedStateUpdate_Done_Inst_n4), .B(Red_RoundConstant[5]), .Z(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_3_n215) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_4_U28 ( 
        .A(Red_RoundConstant[0]), .B(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_4_n71), .ZN(Red_FSMUpdate[4]) );
  AOI22_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_4_U27 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_4_n70), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_4_n69), 
        .B1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_4_n68), .B2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_4_n67), 
        .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_4_n71) );
  OAI21_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_4_U26 ( 
        .B1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_4_n66), .B2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_4_n65), 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_4_n64), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_4_n68)
         );
  AOI21_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_4_U25 ( 
        .B1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_4_n63), .B2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_4_n62), 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_4_n61), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_4_n66)
         );
  AND3_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_4_U24 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_4_n60), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_4_n59), 
        .A3(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_4_n58), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_4_n61)
         );
  OAI21_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_4_U23 ( 
        .B1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_4_n58), .B2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_4_n57), 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_4_n56), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_4_n69)
         );
  NAND3_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_4_U22 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_4_n58), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_4_n55), 
        .A3(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_4_n63), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_4_n56)
         );
  NAND3_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_4_U21 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_4_n62), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_4_n59), 
        .A3(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_4_n67), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_4_n57)
         );
  OAI221_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_4_U20 ( 
        .B1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_4_n54), .B2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_4_n53), 
        .C1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_4_n52), .C2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_4_n51), 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_4_n55), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_4_n67)
         );
  INV_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_4_U19 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_4_n64), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_4_n55)
         );
  XOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_4_U18 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_4_n50), .B(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_4_n49), 
        .Z(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_4_n64) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_4_U17 ( 
        .A(Red_RoundConstant[0]), .B(F_SD2_RedStateUpdate_Done_Inst_n3), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_4_n50) );
  AND2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_4_U16 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_4_n54), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_4_n53), 
        .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_4_n51) );
  OR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_4_U15 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_4_n58), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_4_n62), 
        .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_4_n52) );
  NAND2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_4_U14 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_4_n60), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_4_n65), 
        .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_4_n53) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_4_U13 ( 
        .A(Red_RoundConstant[4]), .B(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_4_n49), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_4_n65)
         );
  XOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_4_U12 ( 
        .A(F_SD2_RedStateUpdate_Done_Inst_n4), .B(
        F_SD2_RedStateUpdate_Done_Inst_n5), .Z(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_4_n49) );
  OR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_4_U11 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_4_n59), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_4_n63), 
        .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_4_n54) );
  XOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_4_U10 ( 
        .A(Red_RoundConstant[6]), .B(F_SD2_RedStateUpdate_Done_Inst_n5), .Z(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_4_n63) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_4_U9 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_4_n48), .B(Red_RoundConstant[1]), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_4_n59) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_4_U8 ( 
        .A(F_SD2_RedStateUpdate_Done_Inst_n3), .B(
        F_SD2_RedStateUpdate_Done_Inst_n4), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_4_n48) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_4_U7 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_4_n47), .B(Red_RoundConstant[2]), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_4_n62) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_4_U6 ( 
        .A(F_SD2_RedStateUpdate_Done_Inst_n3), .B(
        F_SD2_RedStateUpdate_Done_Inst_n5), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_4_n47) );
  XOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_4_U5 ( 
        .A(F_SD2_RedStateUpdate_Done_Inst_n4), .B(Red_RoundConstant[5]), .Z(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_4_n58) );
  INV_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_4_U4 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_4_n60), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_4_n70)
         );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_4_U3 ( 
        .A(F_SD2_RedStateUpdate_Done_Inst_n3), .B(Red_RoundConstant[3]), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_4_n60) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_U56 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n125), .B(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n124), 
        .ZN(Red_FSMUpdate[5]) );
  OAI221_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_U55 ( 
        .B1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n123), .B2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n122), .C1(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n121), .C2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n120), .A(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n119), 
        .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n124) );
  OAI22_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_U54 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n118), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n117), .B1(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n116), .B2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n115), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n119) );
  AND3_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_U53 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n118), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n117), .A3(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n114), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n115) );
  INV_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_U52 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n113), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n116) );
  NOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_U51 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n112), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n111), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n117) );
  AOI21_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_U50 ( 
        .B1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n110), .B2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n109), .A(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n108), 
        .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n122) );
  NOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_U49 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n107), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n106), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n110) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_U48 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n105), .B(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n104), 
        .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n125) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_U47 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n103), .B(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n102), 
        .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n104) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_U46 ( 
        .A(Red_RoundConstant[2]), .B(Red_RoundConstant[5]), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n102) );
  XOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_U45 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n101), .B(Red_RoundConstant[1]), .Z(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n103) );
  AOI211_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_U44 ( 
        .C1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n100), .C2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n99), 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n98), .B(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n97), 
        .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n101) );
  OAI221_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_U43 ( 
        .B1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n96), .B2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n95), 
        .C1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n96), .C2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n94), 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n93), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n97)
         );
  OAI221_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_U42 ( 
        .B1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n92), .B2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n112), .C1(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n92), 
        .C2(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n91), .A(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n96), 
        .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n93) );
  NOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_U41 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n90), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n106), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n92)
         );
  NAND2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_U40 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n111), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n89), 
        .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n106) );
  OR3_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_U39 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n88), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n112), .A3(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n123), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n94)
         );
  INV_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_U38 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n87), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n95)
         );
  NOR3_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_U37 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n86), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n121), .A3(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n113), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n98)
         );
  NAND3_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_U36 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n114), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n88), 
        .A3(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n96), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n113) );
  AOI21_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_U35 ( 
        .B1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n89), .B2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n85), 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n84), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n105) );
  OAI21_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_U34 ( 
        .B1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n83), .B2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n89), 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n82), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n84)
         );
  OAI221_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_U33 ( 
        .B1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n87), .B2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n81), 
        .C1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n87), .C2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n99), 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n112), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n82)
         );
  NAND2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_U32 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n80), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n79), 
        .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n99) );
  INV_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_U31 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n107), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n81)
         );
  NAND2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_U30 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n78), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n96), 
        .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n107) );
  NOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_U29 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n80), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n79), 
        .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n87) );
  NAND2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_U28 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n88), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n86), 
        .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n79) );
  INV_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_U27 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n118), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n80)
         );
  NOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_U26 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n89), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n123), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n118) );
  INV_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_U25 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n121), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n123) );
  AOI21_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_U24 ( 
        .B1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n91), .B2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n100), .A(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n108), 
        .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n83) );
  NOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_U23 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n78), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n90), 
        .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n108) );
  NAND2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_U22 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n112), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n88), 
        .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n90) );
  NOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_U21 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n88), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n121), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n91)
         );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_U20 ( 
        .A(F_SD2_RedStateUpdate_Done_Inst_n3), .B(Red_RoundConstant[3]), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n121) );
  INV_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_U19 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n109), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n88)
         );
  INV_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_U18 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n120), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n85)
         );
  AOI21_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_U17 ( 
        .B1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n100), .B2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n111), .A(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n77), 
        .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n120) );
  AND3_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_U16 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n114), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n109), .A3(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n112), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n77)
         );
  XOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_U15 ( 
        .A(F_SD2_RedStateUpdate_Done_Inst_n5), .B(Red_RoundConstant[6]), .Z(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n109) );
  INV_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_U14 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n86), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n111) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_U13 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n76), .B(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n75), 
        .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n86) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_U12 ( 
        .A(F_SD2_RedStateUpdate_Done_Inst_n5), .B(Red_RoundConstant[0]), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n76) );
  NOR3_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_U11 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n96), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n114), .A3(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n112), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n100) );
  XOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_U10 ( 
        .A(Red_RoundConstant[5]), .B(F_SD2_RedStateUpdate_Done_Inst_n4), .Z(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n112) );
  INV_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_U9 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n78), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n114) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_U8 ( 
        .A(F_SD2_RedStateUpdate_Done_Inst_n3), .B(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n74), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n78)
         );
  XOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_U7 ( 
        .A(Red_RoundConstant[2]), .B(F_SD2_RedStateUpdate_Done_Inst_n5), .Z(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n74) );
  XOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_U6 ( 
        .A(Red_RoundConstant[1]), .B(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n75), .Z(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n96)
         );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_U5 ( 
        .A(F_SD2_RedStateUpdate_Done_Inst_n3), .B(
        F_SD2_RedStateUpdate_Done_Inst_n4), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n75) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_U4 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n73), .B(Red_RoundConstant[4]), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n89) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_U3 ( 
        .A(F_SD2_RedStateUpdate_Done_Inst_n5), .B(
        F_SD2_RedStateUpdate_Done_Inst_n4), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_5_n73) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_U68 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n151), .B(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n150), 
        .ZN(Red_FSMUpdate[6]) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_U67 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n149), .B(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n148), 
        .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n150) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_U66 ( 
        .A(Red_RoundConstant[1]), .B(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n147), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n148) );
  AOI221_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_U65 ( 
        .B1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n146), .B2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n145), .C1(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n144), .C2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n143), .A(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n142), 
        .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n147) );
  NOR3_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_U64 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n141), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n140), .A3(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n139), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n142) );
  NAND3_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_U63 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n138), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n137), .A3(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n136), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n144) );
  NAND3_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_U62 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n141), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n135), .A3(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n134), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n136) );
  NAND2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_U61 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n133), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n132), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n134) );
  AOI22_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_U60 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n131), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n130), .B1(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n129), .B2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n128), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n138) );
  NOR3_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_U59 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n127), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n126), .A3(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n125), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n146) );
  XOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_U58 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n124), .B(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n123), 
        .Z(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n149) );
  AOI22_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_U57 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n122), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n121), .B1(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n120), .B2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n119), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n123) );
  OAI21_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_U56 ( 
        .B1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n118), .B2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n117), .A(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n126), 
        .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n119) );
  OAI221_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_U55 ( 
        .B1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n143), .B2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n116), .C1(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n145), .C2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n115), .A(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n114), 
        .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n121) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_U54 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n113), .B(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n112), 
        .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n115) );
  AOI22_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_U53 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n130), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n111), .B1(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n131), .B2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n141), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n116) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_U52 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n110), .B(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n109), 
        .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n124) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_U51 ( 
        .A(Red_RoundConstant[0]), .B(Red_RoundConstant[5]), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n109) );
  XOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_U50 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n108), .B(Red_RoundConstant[2]), .Z(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n110) );
  AOI211_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_U49 ( 
        .C1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n107), .C2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n106), .A(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n105), 
        .B(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n104), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n108) );
  OAI211_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_U48 ( 
        .C1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n139), .C2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n133), .A(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n103), 
        .B(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n102), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n104) );
  OR3_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_U47 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n135), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n132), .A3(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n126), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n102) );
  NAND2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_U46 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n101), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n118), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n126) );
  AOI22_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_U45 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n100), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n111), .B1(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n120), .B2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n99), 
        .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n103) );
  INV_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_U44 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n139), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n120) );
  NAND2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_U43 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n127), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n98), 
        .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n139) );
  AOI221_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_U42 ( 
        .B1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n122), .B2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n114), .C1(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n125), .C2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n114), .A(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n111), 
        .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n105) );
  INV_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_U41 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n127), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n111) );
  NAND2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_U40 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n113), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n140), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n125) );
  NAND2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_U39 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n130), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n99), 
        .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n114) );
  NOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_U38 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n101), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n113), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n99)
         );
  NOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_U37 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n141), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n132), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n107) );
  OAI221_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_U36 ( 
        .B1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n101), .B2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n97), 
        .C1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n141), .C2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n137), .A(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n96), 
        .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n151) );
  OAI221_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_U35 ( 
        .B1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n130), .B2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n131), .C1(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n98), 
        .C2(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n95), .A(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n101), 
        .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n96) );
  NOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_U34 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n133), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n132), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n95)
         );
  INV_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_U33 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n131), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n132) );
  INV_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_U32 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n130), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n133) );
  NOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_U31 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n122), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n143), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n98)
         );
  NOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_U30 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n113), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n127), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n131) );
  NOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_U29 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n94), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n118), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n130) );
  INV_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_U28 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n100), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n137) );
  NOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_U27 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n135), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n117), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n100) );
  NAND2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_U26 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n113), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n94), 
        .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n117) );
  INV_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_U25 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n128), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n113) );
  AOI22_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_U24 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n127), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n93), 
        .B1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n143), .B2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n92), 
        .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n97) );
  NOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_U23 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n128), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n112), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n92)
         );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_U22 ( 
        .A(F_SD2_RedStateUpdate_Done_Inst_n5), .B(Red_RoundConstant[6]), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n128) );
  INV_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_U21 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n91), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n93)
         );
  AOI22_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_U20 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n135), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n106), .B1(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n129), .B2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n118), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n91)
         );
  INV_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_U19 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n112), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n118) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_U18 ( 
        .A(Red_RoundConstant[4]), .B(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n90), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n112) );
  XOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_U17 ( 
        .A(F_SD2_RedStateUpdate_Done_Inst_n5), .B(
        F_SD2_RedStateUpdate_Done_Inst_n4), .Z(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n90) );
  NOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_U16 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n135), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n94), 
        .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n129) );
  NOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_U15 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n140), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n145), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n106) );
  INV_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_U14 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n143), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n145) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_U13 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n89), .B(Red_RoundConstant[2]), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n143) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_U12 ( 
        .A(F_SD2_RedStateUpdate_Done_Inst_n5), .B(
        F_SD2_RedStateUpdate_Done_Inst_n3), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n89) );
  INV_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_U11 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n94), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n140) );
  XOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_U10 ( 
        .A(F_SD2_RedStateUpdate_Done_Inst_n3), .B(Red_RoundConstant[3]), .Z(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n94) );
  INV_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_U9 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n122), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n135) );
  XOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_U8 ( 
        .A(F_SD2_RedStateUpdate_Done_Inst_n4), .B(Red_RoundConstant[5]), .Z(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n122) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_U7 ( 
        .A(Red_RoundConstant[1]), .B(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n88), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n127) );
  INV_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_U6 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n141), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n101) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_U5 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n87), .B(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n88), 
        .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n141) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_U4 ( 
        .A(F_SD2_RedStateUpdate_Done_Inst_n4), .B(
        F_SD2_RedStateUpdate_Done_Inst_n3), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n88) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_U3 ( 
        .A(Red_RoundConstant[0]), .B(F_SD2_RedStateUpdate_Done_Inst_n5), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_6_n87) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_U49 ( 
        .A(Red_RoundConstant[8]), .B(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n140), .ZN(Red_FSMUpdate[7]) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_U48 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n139), .B(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n138), 
        .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n140) );
  NAND2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_U47 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n137), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n136), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n138) );
  AOI221_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_U46 ( 
        .B1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n135), .B2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n134), .C1(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n133), .C2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n134), .A(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n132), 
        .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n136) );
  NOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_U45 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n131), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n130), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n132) );
  NAND2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_U44 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n129), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n128), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n131) );
  NOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_U43 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n128), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n127), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n133) );
  AND2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_U42 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n126), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n125), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n135) );
  AOI221_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_U41 ( 
        .B1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n124), .B2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n123), .C1(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n122), .C2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n123), .A(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n121), 
        .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n137) );
  NOR4_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_U40 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n120), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n128), .A3(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n119), .A4(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n118), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n121) );
  AOI21_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_U39 ( 
        .B1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n117), .B2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n126), .A(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n125), 
        .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n119) );
  NOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_U38 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n116), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n115), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n125) );
  NOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_U37 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n114), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n126), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n122) );
  AND2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_U36 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n113), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n115), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n123) );
  NOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_U35 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n117), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n112), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n124) );
  XOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_U34 ( 
        .A(Red_RoundConstant[9]), .B(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n111), .Z(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n139)
         );
  OAI21_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_U33 ( 
        .B1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n110), .B2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n126), .A(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n109), 
        .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n111) );
  NAND3_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_U32 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n108), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n115), .A3(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n126), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n109) );
  OAI21_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_U31 ( 
        .B1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n114), .B2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n107), .A(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n106), 
        .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n108) );
  OR3_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_U30 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n128), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n130), .A3(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n112), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n106) );
  NAND2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_U29 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n116), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n118), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n130) );
  INV_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_U28 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n134), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n107) );
  NOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_U27 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n129), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n118), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n134) );
  XOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_U26 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n105), .B(F_SD2_RedStateUpdate_Done_Inst_n6), .Z(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n126) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_U25 ( 
        .A(Red_RoundConstant[9]), .B(F_SD2_RedStateUpdate_Done_Inst_n8), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n105) );
  AOI21_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_U24 ( 
        .B1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n113), .B2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n104), .A(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n103), 
        .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n110) );
  OAI22_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_U23 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n117), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n102), .B1(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n128), .B2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n101), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n103) );
  OAI21_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_U22 ( 
        .B1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n113), .B2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n104), .A(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n112), 
        .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n101) );
  INV_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_U21 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n120), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n112) );
  XOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_U20 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n100), .B(Red_RoundConstant[11]), .Z(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n120) );
  INV_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_U19 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n114), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n128) );
  XOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_U18 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n114), .B(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n127), 
        .Z(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n102) );
  XOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_U17 ( 
        .A(Red_RoundConstant[10]), .B(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n99), .Z(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n114)
         );
  NOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_U16 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n115), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n129), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n104) );
  INV_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_U15 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n117), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n129) );
  XOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_U14 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n98), .B(Red_RoundConstant[12]), .Z(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n117) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_U13 ( 
        .A(F_SD2_RedStateUpdate_Done_Inst_n9), .B(
        F_SD2_RedStateUpdate_Done_Inst_n7), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n98) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_U12 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n97), .B(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n100), 
        .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n115) );
  XOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_U11 ( 
        .A(F_SD2_RedStateUpdate_Done_Inst_n8), .B(
        F_SD2_RedStateUpdate_Done_Inst_n7), .Z(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n100) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_U10 ( 
        .A(F_SD2_RedStateUpdate_Done_Inst_n6), .B(Red_RoundConstant[7]), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n97) );
  AND2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_U9 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n127), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n118), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n113) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_U8 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n96), .B(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n99), 
        .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n118) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_U7 ( 
        .A(F_SD2_RedStateUpdate_Done_Inst_n9), .B(
        F_SD2_RedStateUpdate_Done_Inst_n6), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n99) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_U6 ( 
        .A(Red_RoundConstant[8]), .B(F_SD2_RedStateUpdate_Done_Inst_n7), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n96) );
  INV_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_U5 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n116), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n127) );
  XOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_U4 ( 
        .A(Red_RoundConstant[13]), .B(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n95), .Z(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n116)
         );
  XOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_U3 ( 
        .A(F_SD2_RedStateUpdate_Done_Inst_n9), .B(
        F_SD2_RedStateUpdate_Done_Inst_n8), .Z(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_7_n95) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_8_U29 ( 
        .A(Red_RoundConstant[9]), .B(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_8_n108), .ZN(Red_FSMUpdate[8]) );
  OAI21_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_8_U28 ( 
        .B1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_8_n107), .B2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_8_n106), .A(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_8_n105), 
        .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_8_n108) );
  OAI21_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_8_U27 ( 
        .B1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_8_n104), .B2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_8_n103), .A(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_8_n107), 
        .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_8_n105) );
  OAI221_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_8_U26 ( 
        .B1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_8_n102), .B2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_8_n101), .C1(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_8_n101), .C2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_8_n100), .A(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_8_n99), 
        .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_8_n103) );
  OAI21_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_8_U25 ( 
        .B1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_8_n98), .B2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_8_n100), .A(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_8_n101), 
        .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_8_n99) );
  NOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_8_U24 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_8_n97), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_8_n96), 
        .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_8_n102) );
  OAI21_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_8_U23 ( 
        .B1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_8_n101), .B2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_8_n95), 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_8_n94), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_8_n106) );
  AOI22_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_8_U22 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_8_n97), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_8_n93), 
        .B1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_8_n98), .B2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_8_n92), 
        .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_8_n94) );
  XOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_8_U21 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_8_n97), .B(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_8_n101), 
        .Z(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_8_n92) );
  AND2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_8_U20 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_8_n100), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_8_n91), 
        .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_8_n93) );
  OAI221_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_8_U19 ( 
        .B1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_8_n91), .B2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_8_n97), 
        .C1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_8_n91), .C2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_8_n100), .A(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_8_n96), 
        .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_8_n95) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_8_U18 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_8_n90), .B(Red_RoundConstant[11]), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_8_n96) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_8_U17 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_8_n89), .B(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_8_n88), 
        .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_8_n100) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_8_U16 ( 
        .A(F_SD2_RedStateUpdate_Done_Inst_n7), .B(Red_RoundConstant[8]), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_8_n89) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_8_U15 ( 
        .A(F_SD2_RedStateUpdate_Done_Inst_n9), .B(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_8_n87), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_8_n97)
         );
  XOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_8_U14 ( 
        .A(F_SD2_RedStateUpdate_Done_Inst_n8), .B(Red_RoundConstant[13]), .Z(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_8_n87) );
  NOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_8_U13 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_8_n98), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_8_n86), 
        .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_8_n91) );
  INV_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_8_U12 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_8_n104), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_8_n86)
         );
  XOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_8_U11 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_8_n85), .B(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_8_n90), 
        .Z(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_8_n104) );
  XOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_8_U10 ( 
        .A(F_SD2_RedStateUpdate_Done_Inst_n8), .B(
        F_SD2_RedStateUpdate_Done_Inst_n7), .Z(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_8_n90) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_8_U9 ( 
        .A(F_SD2_RedStateUpdate_Done_Inst_n6), .B(Red_RoundConstant[7]), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_8_n85) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_8_U8 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_8_n84), .B(Red_RoundConstant[12]), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_8_n98) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_8_U7 ( 
        .A(F_SD2_RedStateUpdate_Done_Inst_n9), .B(
        F_SD2_RedStateUpdate_Done_Inst_n7), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_8_n84) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_8_U6 ( 
        .A(Red_RoundConstant[10]), .B(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_8_n88), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_8_n101) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_8_U5 ( 
        .A(F_SD2_RedStateUpdate_Done_Inst_n9), .B(
        F_SD2_RedStateUpdate_Done_Inst_n6), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_8_n88) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_8_U4 ( 
        .A(Red_RoundConstant[9]), .B(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_8_n83), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_8_n107) );
  XOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_8_U3 ( 
        .A(F_SD2_RedStateUpdate_Done_Inst_n8), .B(
        F_SD2_RedStateUpdate_Done_Inst_n6), .Z(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_8_n83) );
  INV_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_9_U33 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_9_n116), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_9_n117) );
  INV_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_9_U32 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_9_n114), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_9_n115) );
  INV_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_9_U31 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_9_n101), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_9_n103) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_9_U30 ( 
        .A(Red_RoundConstant[12]), .B(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_9_n119), .ZN(Red_FSMUpdate[9]) );
  AOI21_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_9_U29 ( 
        .B1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_9_n91), .B2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_9_n109), .A(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_9_n118), 
        .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_9_n119) );
  MUX2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_9_U28 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_9_n112), .B(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_9_n117), 
        .S(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_9_n105), .Z(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_9_n118)
         );
  AOI21_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_9_U27 ( 
        .B1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_9_n104), .B2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_9_n98), 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_9_n115), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_9_n116) );
  OAI211_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_9_U26 ( 
        .C1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_9_n97), .C2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_9_n91), 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_9_n102), .B(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_9_n113), 
        .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_9_n114) );
  OR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_9_U25 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_9_n96), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_9_n109), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_9_n113) );
  NOR3_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_9_U24 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_9_n102), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_9_n111), .A3(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_9_n101), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_9_n112) );
  OAI21_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_9_U23 ( 
        .B1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_9_n94), .B2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_9_n91), 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_9_n110), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_9_n111) );
  OAI21_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_9_U22 ( 
        .B1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_9_n107), .B2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_9_n96), 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_9_n91), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_9_n110) );
  INV_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_9_U21 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_9_n96), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_9_n97)
         );
  NAND2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_9_U20 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_9_n91), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_9_n108), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_9_n109) );
  OAI211_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_9_U19 ( 
        .C1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_9_n98), .C2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_9_n104), .A(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_9_n105), 
        .B(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_9_n107), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_9_n108) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_9_U18 ( 
        .A(F_SD2_RedStateUpdate_Done_Inst_n6), .B(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_9_n106), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_9_n107) );
  XOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_9_U17 ( 
        .A(Red_RoundConstant[10]), .B(F_SD2_RedStateUpdate_Done_Inst_n9), .Z(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_9_n106) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_9_U16 ( 
        .A(Red_RoundConstant[12]), .B(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_9_n99), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_9_n105) );
  NOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_9_U15 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_9_n103), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_9_n102), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_9_n104) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_9_U14 ( 
        .A(Red_RoundConstant[9]), .B(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_9_n92), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_9_n102) );
  XOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_9_U13 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_9_n100), .B(Red_RoundConstant[8]), .Z(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_9_n101) );
  XOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_9_U12 ( 
        .A(F_SD2_RedStateUpdate_Done_Inst_n6), .B(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_9_n99), .Z(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_9_n100)
         );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_9_U11 ( 
        .A(F_SD2_RedStateUpdate_Done_Inst_n7), .B(
        F_SD2_RedStateUpdate_Done_Inst_n9), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_9_n99) );
  NOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_9_U10 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_9_n94), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_9_n97), 
        .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_9_n98) );
  XOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_9_U9 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_9_n95), .B(Red_RoundConstant[13]), .Z(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_9_n96) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_9_U8 ( 
        .A(F_SD2_RedStateUpdate_Done_Inst_n8), .B(
        F_SD2_RedStateUpdate_Done_Inst_n9), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_9_n95) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_9_U7 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_9_n93), .B(Red_RoundConstant[7]), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_9_n94) );
  XOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_9_U6 ( 
        .A(F_SD2_RedStateUpdate_Done_Inst_n7), .B(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_9_n92), .Z(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_9_n93)
         );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_9_U5 ( 
        .A(F_SD2_RedStateUpdate_Done_Inst_n8), .B(
        F_SD2_RedStateUpdate_Done_Inst_n6), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_9_n92) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_9_U4 ( 
        .A(F_SD2_RedStateUpdate_Done_Inst_n8), .B(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_9_n90), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_9_n91)
         );
  XOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_9_U3 ( 
        .A(Red_RoundConstant[11]), .B(F_SD2_RedStateUpdate_Done_Inst_n7), .Z(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_9_n90) );
  INV_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_U47 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n126), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n130) );
  XOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_U46 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n124), .B(F_SD2_RedStateUpdate_Done_Inst_n7), .Z(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n126) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_U45 ( 
        .A(Red_RoundConstant[12]), .B(F_SD2_RedStateUpdate_Done_Inst_n9), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n124) );
  INV_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_U44 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n129), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n127) );
  XOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_U43 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n123), .B(Red_RoundConstant[9]), .Z(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n129) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_U42 ( 
        .A(F_SD2_RedStateUpdate_Done_Inst_n8), .B(
        F_SD2_RedStateUpdate_Done_Inst_n6), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n123) );
  INV_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_U41 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n125), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n128) );
  XOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_U40 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n122), .B(Red_RoundConstant[10]), .Z(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n125) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_U39 ( 
        .A(F_SD2_RedStateUpdate_Done_Inst_n9), .B(
        F_SD2_RedStateUpdate_Done_Inst_n6), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n122) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_U38 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n120), .B(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n121), .ZN(Red_FSMUpdate[10]) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_U37 ( 
        .A(Red_RoundConstant[8]), .B(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n109), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n121) );
  XOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_U36 ( 
        .A(Red_RoundConstant[12]), .B(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n119), .Z(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n120) );
  AOI21_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_U35 ( 
        .B1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n111), .B2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n90), .A(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n118), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n119) );
  OAI21_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_U34 ( 
        .B1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n113), .B2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n90), .A(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n117), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n118) );
  OAI22_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_U33 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n114), .A2(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n115), .B1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n105), .B2(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n116), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n117) );
  AND3_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_U32 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n114), .A2(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n115), .A3(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n97), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n116) );
  NOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_U31 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n101), .A2(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n128), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n115) );
  INV_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_U30 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n94), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n114) );
  OAI221_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_U29 ( 
        .B1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n125), .B2(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n130), .C1(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n97), .C2(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n128), .A(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n112), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n113) );
  NAND2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_U28 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n130), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n97), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n112) );
  AOI211_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_U27 ( 
        .C1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n107), .C2(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n110), .A(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n97), 
        .B(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n93), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n111) );
  NAND2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_U26 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n127), .A2(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n128), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n110) );
  AOI211_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_U25 ( 
        .C1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n130), .C2(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n102), .A(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n104), .B(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n108), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n109) );
  AOI221_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_U24 ( 
        .B1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n129), .B2(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n106), .C1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n107), .C2(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n106), .A(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n90), 
        .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n108) );
  NAND2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_U23 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n101), .A2(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n130), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n107) );
  NAND3_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_U22 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n105), .A2(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n128), .A3(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n88), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n106) );
  INV_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_U21 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n103), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n105) );
  NOR3_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_U20 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n103), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n93), .A3(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n88), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n104) );
  INV_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_U19 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n88), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n101) );
  NAND3_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_U18 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n126), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n97), .A3(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n95), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n103) );
  OAI22_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_U17 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n101), .A2(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n100), .B1(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n98), .B2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n94), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n102) );
  AOI21_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_U16 ( 
        .B1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n127), .B2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n90), .A(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n99), 
        .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n100) );
  AOI21_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_U15 ( 
        .B1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n94), .B2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n98), .A(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n128), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n99) );
  OR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_U14 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n127), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n97), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n98) );
  XOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_U13 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n96), .B(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n91), 
        .Z(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n97) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_U12 ( 
        .A(Red_RoundConstant[8]), .B(F_SD2_RedStateUpdate_Done_Inst_n9), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n96) );
  INV_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_U11 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n127), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n95) );
  NAND2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_U10 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n93), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n90), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n94) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_U9 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n92), .B(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n91), 
        .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n93) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_U8 ( 
        .A(F_SD2_RedStateUpdate_Done_Inst_n8), .B(Red_RoundConstant[7]), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n92) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_U7 ( 
        .A(F_SD2_RedStateUpdate_Done_Inst_n7), .B(
        F_SD2_RedStateUpdate_Done_Inst_n6), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n91) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_U6 ( 
        .A(Red_RoundConstant[13]), .B(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n89), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n90) );
  XOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_U5 ( 
        .A(F_SD2_RedStateUpdate_Done_Inst_n9), .B(
        F_SD2_RedStateUpdate_Done_Inst_n8), .Z(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n89) );
  XOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_U4 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n87), .B(Red_RoundConstant[11]), .Z(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n88) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_U3 ( 
        .A(F_SD2_RedStateUpdate_Done_Inst_n7), .B(
        F_SD2_RedStateUpdate_Done_Inst_n8), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_10_n87) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_U45 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n124), .B(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n123), .ZN(Red_FSMUpdate[11]) );
  OAI211_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_U44 ( 
        .C1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n122), .C2(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n121), .A(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n120), .B(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n119), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n123) );
  OAI22_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_U43 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n118), .A2(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n117), .B1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n116), .B2(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n115), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n119) );
  NOR3_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_U42 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n114), .A2(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n113), .A3(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n121), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n115) );
  INV_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_U41 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n117), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n113) );
  INV_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_U40 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n114), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n118) );
  OAI221_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_U39 ( 
        .B1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n112), .B2(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n111), .C1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n112), .C2(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n110), .A(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n121), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n120) );
  AOI211_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_U38 ( 
        .C1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n109), .C2(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n108), .A(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n117), .B(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n107), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n110) );
  NOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_U37 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n106), .A2(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n105), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n117) );
  INV_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_U36 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n104), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n108) );
  NOR3_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_U35 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n103), .A2(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n102), .A3(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n101), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n112) );
  INV_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_U34 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n105), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n101) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_U33 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n100), .B(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n99), 
        .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n124) );
  AOI21_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_U32 ( 
        .B1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n111), .B2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n98), .A(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n97), 
        .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n99) );
  OAI21_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_U31 ( 
        .B1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n122), .B2(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n111), .A(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n96), 
        .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n97) );
  OAI221_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_U30 ( 
        .B1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n104), .B2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n95), .C1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n104), .C2(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n105), .A(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n116), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n96) );
  NOR3_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_U29 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n94), .A2(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n111), .A3(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n121), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n116) );
  INV_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_U28 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n109), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n95) );
  NOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_U27 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n103), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n93), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n104) );
  NAND2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_U26 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n94), .A2(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n107), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n122) );
  NOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_U25 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n109), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n93), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n107) );
  INV_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_U24 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n106), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n93) );
  OAI22_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_U23 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n106), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n92), .B1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n114), .B2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n91), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n98) );
  AOI21_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_U22 ( 
        .B1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n94), .B2(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n109), .A(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n90), 
        .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n92) );
  AOI21_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_U21 ( 
        .B1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n114), .B2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n91), .A(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n105), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n90) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_U20 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n89), .B(Red_RoundConstant[11]), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n105) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_U19 ( 
        .A(F_SD2_RedStateUpdate_Done_Inst_n7), .B(
        F_SD2_RedStateUpdate_Done_Inst_n8), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n89) );
  NAND2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_U18 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n102), .A2(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n121), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n91) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_U17 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n88), .B(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n87), 
        .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n121) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_U16 ( 
        .A(Red_RoundConstant[7]), .B(F_SD2_RedStateUpdate_Done_Inst_n7), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n88) );
  INV_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_U15 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n94), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n102) );
  NAND2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_U14 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n109), .A2(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n103), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n114) );
  XOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_U13 ( 
        .A(Red_RoundConstant[9]), .B(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n87), .Z(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n103) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_U12 ( 
        .A(F_SD2_RedStateUpdate_Done_Inst_n6), .B(
        F_SD2_RedStateUpdate_Done_Inst_n8), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n87) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_U11 ( 
        .A(Red_RoundConstant[12]), .B(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n86), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n109) );
  XOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_U10 ( 
        .A(F_SD2_RedStateUpdate_Done_Inst_n7), .B(
        F_SD2_RedStateUpdate_Done_Inst_n9), .Z(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n86) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_U9 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n85), .B(Red_RoundConstant[13]), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n94) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_U8 ( 
        .A(F_SD2_RedStateUpdate_Done_Inst_n9), .B(
        F_SD2_RedStateUpdate_Done_Inst_n8), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n85) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_U7 ( 
        .A(Red_RoundConstant[10]), .B(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n84), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n106) );
  XOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_U6 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n83), .B(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n84), 
        .Z(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n111) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_U5 ( 
        .A(F_SD2_RedStateUpdate_Done_Inst_n9), .B(
        F_SD2_RedStateUpdate_Done_Inst_n6), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n84) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_U4 ( 
        .A(Red_RoundConstant[8]), .B(F_SD2_RedStateUpdate_Done_Inst_n7), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n83) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_U3 ( 
        .A(Red_RoundConstant[7]), .B(Red_RoundConstant[8]), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_11_n100) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_12_U31 ( 
        .A(Red_RoundConstant[7]), .B(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_12_n111), .ZN(Red_FSMUpdate[12]) );
  OAI21_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_12_U30 ( 
        .B1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_12_n86), .B2(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_12_n109), .A(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_12_n110), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_12_n111) );
  NAND3_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_12_U29 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_12_n86), .A2(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_12_n105), .A3(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_12_n95), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_12_n110) );
  OAI21_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_12_U28 ( 
        .B1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_12_n107), .B2(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_12_n101), .A(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_12_n108), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_12_n109) );
  NAND4_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_12_U27 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_12_n94), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_12_n98), .A3(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_12_n96), .A4(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_12_n90), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_12_n108) );
  AOI21_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_12_U26 ( 
        .B1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_12_n96), .B2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_12_n88), .A(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_12_n106), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_12_n107) );
  AND3_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_12_U25 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_12_n92), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_12_n93), .A3(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_12_n98), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_12_n106) );
  INV_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_12_U24 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_12_n90), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_12_n93) );
  NAND2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_12_U23 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_12_n103), .A2(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_12_n104), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_12_n105) );
  OAI22_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_12_U22 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_12_n102), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_12_n99), .B1(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_12_n93), .B2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_12_n96), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_12_n104) );
  NAND2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_12_U21 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_12_n102), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_12_n99), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_12_n103) );
  NAND2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_12_U20 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_12_n92), .A2(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_12_n101), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_12_n102) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_12_U19 ( 
        .A(Red_RoundConstant[9]), .B(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_12_n100), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_12_n101) );
  XOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_12_U18 ( 
        .A(F_SD2_RedStateUpdate_Done_Inst_n8), .B(
        F_SD2_RedStateUpdate_Done_Inst_n6), .Z(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_12_n100) );
  INV_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_12_U17 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_12_n92), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_12_n94) );
  OR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_12_U16 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_12_n88), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_12_n98), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_12_n99) );
  XOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_12_U15 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_12_n97), .B(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_12_n91), 
        .Z(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_12_n98) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_12_U14 ( 
        .A(F_SD2_RedStateUpdate_Done_Inst_n6), .B(Red_RoundConstant[8]), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_12_n97) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_12_U13 ( 
        .A(Red_RoundConstant[11]), .B(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_12_n84), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_12_n96) );
  NAND3_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_12_U12 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_12_n88), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_12_n93), .A3(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_12_n94), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_12_n95) );
  XOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_12_U11 ( 
        .A(Red_RoundConstant[12]), .B(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_12_n91), .Z(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_12_n92)
         );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_12_U10 ( 
        .A(F_SD2_RedStateUpdate_Done_Inst_n9), .B(
        F_SD2_RedStateUpdate_Done_Inst_n7), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_12_n91) );
  XOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_12_U9 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_12_n89), .B(F_SD2_RedStateUpdate_Done_Inst_n6), .Z(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_12_n90) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_12_U8 ( 
        .A(F_SD2_RedStateUpdate_Done_Inst_n9), .B(Red_RoundConstant[10]), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_12_n89) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_12_U7 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_12_n87), .B(Red_RoundConstant[13]), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_12_n88) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_12_U6 ( 
        .A(F_SD2_RedStateUpdate_Done_Inst_n8), .B(
        F_SD2_RedStateUpdate_Done_Inst_n9), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_12_n87) );
  XOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_12_U5 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_12_n85), .B(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_12_n84), 
        .Z(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_12_n86) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_12_U4 ( 
        .A(Red_RoundConstant[7]), .B(F_SD2_RedStateUpdate_Done_Inst_n6), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_12_n85) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_12_U3 ( 
        .A(F_SD2_RedStateUpdate_Done_Inst_n8), .B(
        F_SD2_RedStateUpdate_Done_Inst_n7), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_12_n84) );
  INV_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_13_U29 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_13_n85), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_13_n86) );
  INV_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_13_U28 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_13_n76), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_13_n79) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_13_U27 ( 
        .A(Red_RoundConstant[8]), .B(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_13_n96), .ZN(Red_FSMUpdate[13]) );
  MUX2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_13_U26 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_13_n88), .B(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_13_n93), 
        .S(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_13_n95), .Z(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_13_n96)
         );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_13_U25 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_13_n94), .B(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_13_n75), 
        .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_13_n95) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_13_U24 ( 
        .A(Red_RoundConstant[8]), .B(F_SD2_RedStateUpdate_Done_Inst_n7), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_13_n94) );
  AOI22_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_13_U23 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_13_n89), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_13_n90), .B1(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_13_n72), .B2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_13_n92), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_13_n93) );
  OAI21_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_13_U22 ( 
        .B1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_13_n76), .B2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_13_n85), .A(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_13_n91), 
        .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_13_n92) );
  OAI21_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_13_U21 ( 
        .B1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_13_n90), .B2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_13_n89), .A(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_13_n78), 
        .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_13_n91) );
  AND2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_13_U20 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_13_n79), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_13_n74), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_13_n90) );
  NOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_13_U19 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_13_n86), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_13_n82), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_13_n89) );
  OAI21_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_13_U18 ( 
        .B1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_13_n83), .B2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_13_n86), .A(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_13_n87), 
        .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_13_n88) );
  OAI21_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_13_U17 ( 
        .B1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_13_n72), .B2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_13_n79), .A(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_13_n86), 
        .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_13_n87) );
  XOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_13_U16 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_13_n84), .B(Red_RoundConstant[13]), .Z(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_13_n85) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_13_U15 ( 
        .A(F_SD2_RedStateUpdate_Done_Inst_n9), .B(
        F_SD2_RedStateUpdate_Done_Inst_n8), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_13_n84) );
  AND2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_13_U14 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_13_n80), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_13_n82), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_13_n83) );
  XOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_13_U13 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_13_n81), .B(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_13_n73), 
        .Z(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_13_n82) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_13_U12 ( 
        .A(F_SD2_RedStateUpdate_Done_Inst_n6), .B(Red_RoundConstant[7]), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_13_n81) );
  OAI22_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_13_U11 ( 
        .A1(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_13_n72), .A2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_13_n74), .B1(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_13_n79), .B2(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_13_n78), .ZN(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_13_n80) );
  XOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_13_U10 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_13_n77), .B(Red_RoundConstant[9]), .Z(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_13_n78) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_13_U9 ( 
        .A(F_SD2_RedStateUpdate_Done_Inst_n8), .B(
        F_SD2_RedStateUpdate_Done_Inst_n6), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_13_n77) );
  XOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_13_U8 ( 
        .A(Red_RoundConstant[10]), .B(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_13_n75), .Z(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_13_n76)
         );
  XOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_13_U7 ( 
        .A(F_SD2_RedStateUpdate_Done_Inst_n9), .B(
        F_SD2_RedStateUpdate_Done_Inst_n6), .Z(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_13_n75) );
  XOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_13_U6 ( 
        .A(Red_RoundConstant[11]), .B(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_13_n73), .Z(F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_13_n74)
         );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_13_U5 ( 
        .A(F_SD2_RedStateUpdate_Done_Inst_n7), .B(
        F_SD2_RedStateUpdate_Done_Inst_n8), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_13_n73) );
  XOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_13_U4 ( 
        .A(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_13_n71), .B(F_SD2_RedStateUpdate_Done_Inst_n7), .Z(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_13_n72) );
  XNOR2_X1 F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_13_U3 ( 
        .A(F_SD2_RedStateUpdate_Done_Inst_n9), .B(Red_RoundConstant[12]), .ZN(
        F_SD2_RedStateUpdate_Done_Inst_F_SD2_RedStateUpdate_Done_bit_inst_13_n71) );
  DFF_X1 Red_FSMRegInst_s_current_state_reg_0_ ( .D(Red_FSMUpdate[0]), .CK(clk), .Q(Red_FSMReg[0]), .QN() );
  DFF_X1 Red_FSMRegInst_s_current_state_reg_1_ ( .D(Red_FSMUpdate[1]), .CK(clk), .Q(Red_FSMReg[1]), .QN() );
  DFF_X1 Red_FSMRegInst_s_current_state_reg_2_ ( .D(Red_FSMUpdate[2]), .CK(clk), .Q(Red_FSMReg[2]), .QN() );
  DFF_X1 Red_FSMRegInst_s_current_state_reg_3_ ( .D(Red_FSMUpdate[3]), .CK(clk), .Q(Red_FSMReg[3]), .QN() );
  DFF_X1 Red_FSMRegInst_s_current_state_reg_4_ ( .D(Red_FSMUpdate[4]), .CK(clk), .Q(Red_FSMReg[4]), .QN() );
  DFF_X1 Red_FSMRegInst_s_current_state_reg_5_ ( .D(Red_FSMUpdate[5]), .CK(clk), .Q(Red_FSMReg[5]), .QN() );
  DFF_X1 Red_FSMRegInst_s_current_state_reg_6_ ( .D(Red_FSMUpdate[6]), .CK(clk), .Q(Red_FSMReg[6]), .QN() );
  DFF_X1 Red_FSMRegInst_s_current_state_reg_7_ ( .D(Red_FSMUpdate[7]), .CK(clk), .Q(Red_FSMReg[7]), .QN() );
  DFF_X1 Red_FSMRegInst_s_current_state_reg_8_ ( .D(Red_FSMUpdate[8]), .CK(clk), .Q(Red_FSMReg[8]), .QN() );
  DFF_X1 Red_FSMRegInst_s_current_state_reg_9_ ( .D(Red_FSMUpdate[9]), .CK(clk), .Q(Red_FSMReg[9]), .QN() );
  DFF_X1 Red_FSMRegInst_s_current_state_reg_10_ ( .D(Red_FSMUpdate[10]), .CK(
        clk), .Q(Red_FSMReg[10]), .QN() );
  DFF_X1 Red_FSMRegInst_s_current_state_reg_11_ ( .D(Red_FSMUpdate[11]), .CK(
        clk), .Q(Red_FSMReg[11]), .QN() );
  DFF_X1 Red_FSMRegInst_s_current_state_reg_12_ ( .D(Red_FSMUpdate[12]), .CK(
        clk), .Q(Red_FSMReg[12]), .QN() );
  DFF_X1 Red_FSMRegInst_s_current_state_reg_13_ ( .D(Red_FSMUpdate[13]), .CK(
        clk), .Q(Red_FSMReg[13]), .QN() );
  NOR2_X1 Red_selectsMUX_MUXInst_0_U2 ( .A1(rst), .A2(
        Red_selectsMUX_MUXInst_0_n4), .ZN(KeyMux_sel_input[0]) );
  INV_X1 Red_selectsMUX_MUXInst_0_U1 ( .A(Red_selectsReg[0]), .ZN(
        Red_selectsMUX_MUXInst_0_n4) );
  NOR2_X1 Red_selectsMUX_MUXInst_1_U2 ( .A1(rst), .A2(
        Red_selectsMUX_MUXInst_1_n4), .ZN(KeyMux_sel_input[1]) );
  INV_X1 Red_selectsMUX_MUXInst_1_U1 ( .A(Red_selectsReg[1]), .ZN(
        Red_selectsMUX_MUXInst_1_n4) );
  NOR2_X1 Red_selectsMUX_MUXInst_2_U3 ( .A1(rst), .A2(
        Red_selectsMUX_MUXInst_2_n5), .ZN(Red_selectsMUX_MUXInst_2_n6) );
  INV_X1 Red_selectsMUX_MUXInst_2_U2 ( .A(Red_selectsReg[2]), .ZN(
        Red_selectsMUX_MUXInst_2_n5) );
  BUF_X2 Red_selectsMUX_MUXInst_2_U1 ( .A(Red_selectsMUX_MUXInst_2_n6), .Z(n3)
         );
  INV_X1 Red_selectsMUX_MUXInst_3_U2 ( .A(Red_selectsReg[3]), .ZN(
        Red_selectsMUX_MUXInst_3_n4) );
  NOR2_X2 Red_selectsMUX_MUXInst_3_U1 ( .A1(rst), .A2(
        Red_selectsMUX_MUXInst_3_n4), .ZN(n4) );
  OAI221_X1 F_SD2_Red_SelectsUpdate_Inst_F_SD2_Red_SelectsUpdate_Bit_Inst_0_U10 ( 
        .B1(
        F_SD2_Red_SelectsUpdate_Inst_F_SD2_Red_SelectsUpdate_Bit_Inst_0_n11), 
        .B2(n5), .C1(
        F_SD2_Red_SelectsUpdate_Inst_F_SD2_Red_SelectsUpdate_Bit_Inst_0_n11), 
        .C2(n3), .A(
        F_SD2_Red_SelectsUpdate_Inst_F_SD2_Red_SelectsUpdate_Bit_Inst_0_n12), 
        .ZN(Red_selectsNext[0]) );
  OR3_X1 F_SD2_Red_SelectsUpdate_Inst_F_SD2_Red_SelectsUpdate_Bit_Inst_0_U9 ( 
        .A1(n7), .A2(n4), .A3(n6), .ZN(
        F_SD2_Red_SelectsUpdate_Inst_F_SD2_Red_SelectsUpdate_Bit_Inst_0_n12)
         );
  AOI211_X1 F_SD2_Red_SelectsUpdate_Inst_F_SD2_Red_SelectsUpdate_Bit_Inst_0_U8 ( 
        .C1(F_SD2_Red_SelectsUpdate_Inst_F_SD2_Red_SelectsUpdate_Bit_Inst_0_n6), .C2(F_SD2_Red_SelectsUpdate_Inst_F_SD2_Red_SelectsUpdate_Bit_Inst_0_n7), .A(
        F_SD2_Red_SelectsUpdate_Inst_F_SD2_Red_SelectsUpdate_Bit_Inst_0_n9), 
        .B(F_SD2_Red_SelectsUpdate_Inst_F_SD2_Red_SelectsUpdate_Bit_Inst_0_n10), .ZN(F_SD2_Red_SelectsUpdate_Inst_F_SD2_Red_SelectsUpdate_Bit_Inst_0_n11) );
  NOR2_X1 F_SD2_Red_SelectsUpdate_Inst_F_SD2_Red_SelectsUpdate_Bit_Inst_0_U7 ( 
        .A1(n4), .A2(n6), .ZN(
        F_SD2_Red_SelectsUpdate_Inst_F_SD2_Red_SelectsUpdate_Bit_Inst_0_n10)
         );
  AOI211_X1 F_SD2_Red_SelectsUpdate_Inst_F_SD2_Red_SelectsUpdate_Bit_Inst_0_U6 ( 
        .C1(F_SD2_Red_SelectsUpdate_Inst_F_SD2_Red_SelectsUpdate_Bit_Inst_0_n8), .C2(n7), .A(n5), .B(n3), .ZN(
        F_SD2_Red_SelectsUpdate_Inst_F_SD2_Red_SelectsUpdate_Bit_Inst_0_n9) );
  INV_X1 F_SD2_Red_SelectsUpdate_Inst_F_SD2_Red_SelectsUpdate_Bit_Inst_0_U5 ( 
        .A(F_SD2_Red_SelectsUpdate_Inst_F_SD2_Red_SelectsUpdate_Bit_Inst_0_n7), 
        .ZN(F_SD2_Red_SelectsUpdate_Inst_F_SD2_Red_SelectsUpdate_Bit_Inst_0_n8) );
  NAND2_X1 F_SD2_Red_SelectsUpdate_Inst_F_SD2_Red_SelectsUpdate_Bit_Inst_0_U4 ( 
        .A1(n4), .A2(n6), .ZN(
        F_SD2_Red_SelectsUpdate_Inst_F_SD2_Red_SelectsUpdate_Bit_Inst_0_n7) );
  INV_X1 F_SD2_Red_SelectsUpdate_Inst_F_SD2_Red_SelectsUpdate_Bit_Inst_0_U3 ( 
        .A(n7), .ZN(
        F_SD2_Red_SelectsUpdate_Inst_F_SD2_Red_SelectsUpdate_Bit_Inst_0_n6) );
  OAI221_X1 F_SD2_Red_SelectsUpdate_Inst_F_SD2_Red_SelectsUpdate_Bit_Inst_1_U10 ( 
        .B1(
        F_SD2_Red_SelectsUpdate_Inst_F_SD2_Red_SelectsUpdate_Bit_Inst_1_n11), 
        .B2(n5), .C1(
        F_SD2_Red_SelectsUpdate_Inst_F_SD2_Red_SelectsUpdate_Bit_Inst_1_n11), 
        .C2(n3), .A(
        F_SD2_Red_SelectsUpdate_Inst_F_SD2_Red_SelectsUpdate_Bit_Inst_1_n12), 
        .ZN(Red_selectsNext[1]) );
  OR3_X1 F_SD2_Red_SelectsUpdate_Inst_F_SD2_Red_SelectsUpdate_Bit_Inst_1_U9 ( 
        .A1(n7), .A2(n4), .A3(n6), .ZN(
        F_SD2_Red_SelectsUpdate_Inst_F_SD2_Red_SelectsUpdate_Bit_Inst_1_n12)
         );
  AOI211_X1 F_SD2_Red_SelectsUpdate_Inst_F_SD2_Red_SelectsUpdate_Bit_Inst_1_U8 ( 
        .C1(F_SD2_Red_SelectsUpdate_Inst_F_SD2_Red_SelectsUpdate_Bit_Inst_1_n6), .C2(F_SD2_Red_SelectsUpdate_Inst_F_SD2_Red_SelectsUpdate_Bit_Inst_1_n7), .A(
        F_SD2_Red_SelectsUpdate_Inst_F_SD2_Red_SelectsUpdate_Bit_Inst_1_n9), 
        .B(F_SD2_Red_SelectsUpdate_Inst_F_SD2_Red_SelectsUpdate_Bit_Inst_1_n10), .ZN(F_SD2_Red_SelectsUpdate_Inst_F_SD2_Red_SelectsUpdate_Bit_Inst_1_n11) );
  NOR2_X1 F_SD2_Red_SelectsUpdate_Inst_F_SD2_Red_SelectsUpdate_Bit_Inst_1_U7 ( 
        .A1(n4), .A2(n6), .ZN(
        F_SD2_Red_SelectsUpdate_Inst_F_SD2_Red_SelectsUpdate_Bit_Inst_1_n10)
         );
  AOI211_X1 F_SD2_Red_SelectsUpdate_Inst_F_SD2_Red_SelectsUpdate_Bit_Inst_1_U6 ( 
        .C1(F_SD2_Red_SelectsUpdate_Inst_F_SD2_Red_SelectsUpdate_Bit_Inst_1_n8), .C2(n7), .A(n5), .B(n3), .ZN(
        F_SD2_Red_SelectsUpdate_Inst_F_SD2_Red_SelectsUpdate_Bit_Inst_1_n9) );
  INV_X1 F_SD2_Red_SelectsUpdate_Inst_F_SD2_Red_SelectsUpdate_Bit_Inst_1_U5 ( 
        .A(F_SD2_Red_SelectsUpdate_Inst_F_SD2_Red_SelectsUpdate_Bit_Inst_1_n7), 
        .ZN(F_SD2_Red_SelectsUpdate_Inst_F_SD2_Red_SelectsUpdate_Bit_Inst_1_n8) );
  NAND2_X1 F_SD2_Red_SelectsUpdate_Inst_F_SD2_Red_SelectsUpdate_Bit_Inst_1_U4 ( 
        .A1(n4), .A2(n6), .ZN(
        F_SD2_Red_SelectsUpdate_Inst_F_SD2_Red_SelectsUpdate_Bit_Inst_1_n7) );
  INV_X1 F_SD2_Red_SelectsUpdate_Inst_F_SD2_Red_SelectsUpdate_Bit_Inst_1_U3 ( 
        .A(n7), .ZN(
        F_SD2_Red_SelectsUpdate_Inst_F_SD2_Red_SelectsUpdate_Bit_Inst_1_n6) );
  OAI221_X1 F_SD2_Red_SelectsUpdate_Inst_F_SD2_Red_SelectsUpdate_Bit_Inst_2_U10 ( 
        .B1(
        F_SD2_Red_SelectsUpdate_Inst_F_SD2_Red_SelectsUpdate_Bit_Inst_2_n28), 
        .B2(n5), .C1(
        F_SD2_Red_SelectsUpdate_Inst_F_SD2_Red_SelectsUpdate_Bit_Inst_2_n28), 
        .C2(n3), .A(
        F_SD2_Red_SelectsUpdate_Inst_F_SD2_Red_SelectsUpdate_Bit_Inst_2_n29), 
        .ZN(Red_selectsNext[2]) );
  OR3_X1 F_SD2_Red_SelectsUpdate_Inst_F_SD2_Red_SelectsUpdate_Bit_Inst_2_U9 ( 
        .A1(n7), .A2(n4), .A3(n6), .ZN(
        F_SD2_Red_SelectsUpdate_Inst_F_SD2_Red_SelectsUpdate_Bit_Inst_2_n29)
         );
  AOI211_X1 F_SD2_Red_SelectsUpdate_Inst_F_SD2_Red_SelectsUpdate_Bit_Inst_2_U8 ( 
        .C1(
        F_SD2_Red_SelectsUpdate_Inst_F_SD2_Red_SelectsUpdate_Bit_Inst_2_n23), 
        .C2(
        F_SD2_Red_SelectsUpdate_Inst_F_SD2_Red_SelectsUpdate_Bit_Inst_2_n24), 
        .A(F_SD2_Red_SelectsUpdate_Inst_F_SD2_Red_SelectsUpdate_Bit_Inst_2_n26), .B(F_SD2_Red_SelectsUpdate_Inst_F_SD2_Red_SelectsUpdate_Bit_Inst_2_n27), 
        .ZN(
        F_SD2_Red_SelectsUpdate_Inst_F_SD2_Red_SelectsUpdate_Bit_Inst_2_n28)
         );
  NOR2_X1 F_SD2_Red_SelectsUpdate_Inst_F_SD2_Red_SelectsUpdate_Bit_Inst_2_U7 ( 
        .A1(n4), .A2(n6), .ZN(
        F_SD2_Red_SelectsUpdate_Inst_F_SD2_Red_SelectsUpdate_Bit_Inst_2_n27)
         );
  AOI211_X1 F_SD2_Red_SelectsUpdate_Inst_F_SD2_Red_SelectsUpdate_Bit_Inst_2_U6 ( 
        .C1(
        F_SD2_Red_SelectsUpdate_Inst_F_SD2_Red_SelectsUpdate_Bit_Inst_2_n25), 
        .C2(n7), .A(n5), .B(n3), .ZN(
        F_SD2_Red_SelectsUpdate_Inst_F_SD2_Red_SelectsUpdate_Bit_Inst_2_n26)
         );
  INV_X1 F_SD2_Red_SelectsUpdate_Inst_F_SD2_Red_SelectsUpdate_Bit_Inst_2_U5 ( 
        .A(F_SD2_Red_SelectsUpdate_Inst_F_SD2_Red_SelectsUpdate_Bit_Inst_2_n24), .ZN(F_SD2_Red_SelectsUpdate_Inst_F_SD2_Red_SelectsUpdate_Bit_Inst_2_n25) );
  NAND2_X1 F_SD2_Red_SelectsUpdate_Inst_F_SD2_Red_SelectsUpdate_Bit_Inst_2_U4 ( 
        .A1(n4), .A2(n6), .ZN(
        F_SD2_Red_SelectsUpdate_Inst_F_SD2_Red_SelectsUpdate_Bit_Inst_2_n24)
         );
  INV_X1 F_SD2_Red_SelectsUpdate_Inst_F_SD2_Red_SelectsUpdate_Bit_Inst_2_U3 ( 
        .A(n7), .ZN(
        F_SD2_Red_SelectsUpdate_Inst_F_SD2_Red_SelectsUpdate_Bit_Inst_2_n23)
         );
  OAI221_X1 F_SD2_Red_SelectsUpdate_Inst_F_SD2_Red_SelectsUpdate_Bit_Inst_3_U10 ( 
        .B1(
        F_SD2_Red_SelectsUpdate_Inst_F_SD2_Red_SelectsUpdate_Bit_Inst_3_n11), 
        .B2(n5), .C1(
        F_SD2_Red_SelectsUpdate_Inst_F_SD2_Red_SelectsUpdate_Bit_Inst_3_n11), 
        .C2(n3), .A(
        F_SD2_Red_SelectsUpdate_Inst_F_SD2_Red_SelectsUpdate_Bit_Inst_3_n12), 
        .ZN(Red_selectsNext[3]) );
  OR3_X1 F_SD2_Red_SelectsUpdate_Inst_F_SD2_Red_SelectsUpdate_Bit_Inst_3_U9 ( 
        .A1(n7), .A2(n4), .A3(n6), .ZN(
        F_SD2_Red_SelectsUpdate_Inst_F_SD2_Red_SelectsUpdate_Bit_Inst_3_n12)
         );
  AOI211_X1 F_SD2_Red_SelectsUpdate_Inst_F_SD2_Red_SelectsUpdate_Bit_Inst_3_U8 ( 
        .C1(F_SD2_Red_SelectsUpdate_Inst_F_SD2_Red_SelectsUpdate_Bit_Inst_3_n6), .C2(F_SD2_Red_SelectsUpdate_Inst_F_SD2_Red_SelectsUpdate_Bit_Inst_3_n7), .A(
        F_SD2_Red_SelectsUpdate_Inst_F_SD2_Red_SelectsUpdate_Bit_Inst_3_n9), 
        .B(F_SD2_Red_SelectsUpdate_Inst_F_SD2_Red_SelectsUpdate_Bit_Inst_3_n10), .ZN(F_SD2_Red_SelectsUpdate_Inst_F_SD2_Red_SelectsUpdate_Bit_Inst_3_n11) );
  NOR2_X1 F_SD2_Red_SelectsUpdate_Inst_F_SD2_Red_SelectsUpdate_Bit_Inst_3_U7 ( 
        .A1(n4), .A2(n6), .ZN(
        F_SD2_Red_SelectsUpdate_Inst_F_SD2_Red_SelectsUpdate_Bit_Inst_3_n10)
         );
  AOI211_X1 F_SD2_Red_SelectsUpdate_Inst_F_SD2_Red_SelectsUpdate_Bit_Inst_3_U6 ( 
        .C1(F_SD2_Red_SelectsUpdate_Inst_F_SD2_Red_SelectsUpdate_Bit_Inst_3_n8), .C2(n7), .A(n5), .B(n3), .ZN(
        F_SD2_Red_SelectsUpdate_Inst_F_SD2_Red_SelectsUpdate_Bit_Inst_3_n9) );
  INV_X1 F_SD2_Red_SelectsUpdate_Inst_F_SD2_Red_SelectsUpdate_Bit_Inst_3_U5 ( 
        .A(F_SD2_Red_SelectsUpdate_Inst_F_SD2_Red_SelectsUpdate_Bit_Inst_3_n7), 
        .ZN(F_SD2_Red_SelectsUpdate_Inst_F_SD2_Red_SelectsUpdate_Bit_Inst_3_n8) );
  NAND2_X1 F_SD2_Red_SelectsUpdate_Inst_F_SD2_Red_SelectsUpdate_Bit_Inst_3_U4 ( 
        .A1(n4), .A2(n6), .ZN(
        F_SD2_Red_SelectsUpdate_Inst_F_SD2_Red_SelectsUpdate_Bit_Inst_3_n7) );
  INV_X1 F_SD2_Red_SelectsUpdate_Inst_F_SD2_Red_SelectsUpdate_Bit_Inst_3_U3 ( 
        .A(n7), .ZN(
        F_SD2_Red_SelectsUpdate_Inst_F_SD2_Red_SelectsUpdate_Bit_Inst_3_n6) );
  DFF_X1 Red_selectsRegInst_s_current_state_reg_0_ ( .D(Red_selectsNext[0]), 
        .CK(clk), .Q(Red_selectsReg[0]), .QN() );
  DFF_X1 Red_selectsRegInst_s_current_state_reg_1_ ( .D(Red_selectsNext[1]), 
        .CK(clk), .Q(Red_selectsReg[1]), .QN() );
  DFF_X1 Red_selectsRegInst_s_current_state_reg_2_ ( .D(Red_selectsNext[2]), 
        .CK(clk), .Q(Red_selectsReg[2]), .QN() );
  DFF_X1 Red_selectsRegInst_s_current_state_reg_3_ ( .D(Red_selectsNext[3]), 
        .CK(clk), .Q(Red_selectsReg[3]), .QN() );
  BUF_X1 Output_MUX_U4 ( .A(Red_done[0]), .Z(Output_MUX_n8) );
  BUF_X1 Output_MUX_U3 ( .A(done), .Z(Output_MUX_n10) );
  BUF_X1 Output_MUX_U2 ( .A(Red_done[0]), .Z(Output_MUX_n7) );
  CLKBUF_X2 Output_MUX_U1 ( .A(Red_done[1]), .Z(Output_MUX_n9) );
  AND4_X1 Output_MUX_AND3_inst_0_U1 ( .A1(Red_done[1]), .A2(OutputRegIn[0]), 
        .A3(Output_MUX_n8), .A4(done), .ZN(Output[0]) );
  AND4_X1 Output_MUX_AND3_inst_1_U1 ( .A1(Output_MUX_n9), .A2(OutputRegIn[1]), 
        .A3(Output_MUX_n7), .A4(done), .ZN(Output[1]) );
  AND4_X1 Output_MUX_AND3_inst_2_U1 ( .A1(Output_MUX_n9), .A2(OutputRegIn[2]), 
        .A3(Output_MUX_n7), .A4(done), .ZN(Output[2]) );
  AND4_X1 Output_MUX_AND3_inst_3_U1 ( .A1(Output_MUX_n9), .A2(OutputRegIn[3]), 
        .A3(Output_MUX_n8), .A4(done), .ZN(Output[3]) );
  AND4_X1 Output_MUX_AND3_inst_4_U1 ( .A1(Output_MUX_n9), .A2(OutputRegIn[4]), 
        .A3(Output_MUX_n7), .A4(Output_MUX_n10), .ZN(Output[4]) );
  AND4_X1 Output_MUX_AND3_inst_5_U1 ( .A1(Output_MUX_n9), .A2(OutputRegIn[5]), 
        .A3(Output_MUX_n8), .A4(done), .ZN(Output[5]) );
  AND4_X1 Output_MUX_AND3_inst_6_U1 ( .A1(Output_MUX_n9), .A2(OutputRegIn[6]), 
        .A3(Output_MUX_n8), .A4(done), .ZN(Output[6]) );
  AND4_X1 Output_MUX_AND3_inst_7_U1 ( .A1(Output_MUX_n9), .A2(OutputRegIn[7]), 
        .A3(Output_MUX_n7), .A4(done), .ZN(Output[7]) );
  AND4_X1 Output_MUX_AND3_inst_8_U1 ( .A1(Output_MUX_n9), .A2(OutputRegIn[8]), 
        .A3(Red_done[0]), .A4(done), .ZN(Output[8]) );
  AND4_X1 Output_MUX_AND3_inst_9_U1 ( .A1(Output_MUX_n9), .A2(OutputRegIn[9]), 
        .A3(Output_MUX_n7), .A4(Output_MUX_n10), .ZN(Output[9]) );
  AND4_X1 Output_MUX_AND3_inst_10_U1 ( .A1(Output_MUX_n9), .A2(OutputRegIn[10]), .A3(Output_MUX_n8), .A4(done), .ZN(Output[10]) );
  AND4_X1 Output_MUX_AND3_inst_11_U1 ( .A1(Output_MUX_n9), .A2(OutputRegIn[11]), .A3(Output_MUX_n7), .A4(done), .ZN(Output[11]) );
  AND4_X1 Output_MUX_AND3_inst_12_U1 ( .A1(Output_MUX_n9), .A2(OutputRegIn[12]), .A3(Red_done[0]), .A4(done), .ZN(Output[12]) );
  AND4_X1 Output_MUX_AND3_inst_13_U1 ( .A1(Output_MUX_n9), .A2(OutputRegIn[13]), .A3(Red_done[0]), .A4(done), .ZN(Output[13]) );
  AND4_X1 Output_MUX_AND3_inst_14_U1 ( .A1(Output_MUX_n9), .A2(OutputRegIn[14]), .A3(Output_MUX_n8), .A4(done), .ZN(Output[14]) );
  AND4_X1 Output_MUX_AND3_inst_15_U1 ( .A1(Output_MUX_n9), .A2(OutputRegIn[15]), .A3(Output_MUX_n8), .A4(done), .ZN(Output[15]) );
  AND4_X1 Output_MUX_AND3_inst_16_U1 ( .A1(Output_MUX_n9), .A2(OutputRegIn[16]), .A3(Output_MUX_n7), .A4(done), .ZN(Output[16]) );
  AND4_X1 Output_MUX_AND3_inst_17_U1 ( .A1(Output_MUX_n9), .A2(OutputRegIn[17]), .A3(Red_done[0]), .A4(done), .ZN(Output[17]) );
  AND4_X1 Output_MUX_AND3_inst_18_U1 ( .A1(Output_MUX_n9), .A2(OutputRegIn[18]), .A3(Red_done[0]), .A4(done), .ZN(Output[18]) );
  AND4_X1 Output_MUX_AND3_inst_19_U1 ( .A1(Output_MUX_n9), .A2(OutputRegIn[19]), .A3(Red_done[0]), .A4(done), .ZN(Output[19]) );
  AND4_X1 Output_MUX_AND3_inst_20_U1 ( .A1(Output_MUX_n9), .A2(OutputRegIn[20]), .A3(Output_MUX_n8), .A4(done), .ZN(Output[20]) );
  AND4_X1 Output_MUX_AND3_inst_21_U1 ( .A1(Output_MUX_n9), .A2(OutputRegIn[21]), .A3(Output_MUX_n7), .A4(done), .ZN(Output[21]) );
  AND4_X1 Output_MUX_AND3_inst_22_U1 ( .A1(Output_MUX_n9), .A2(OutputRegIn[22]), .A3(Red_done[0]), .A4(done), .ZN(Output[22]) );
  AND4_X1 Output_MUX_AND3_inst_23_U1 ( .A1(Output_MUX_n9), .A2(OutputRegIn[23]), .A3(Red_done[0]), .A4(done), .ZN(Output[23]) );
  AND4_X1 Output_MUX_AND3_inst_24_U1 ( .A1(Output_MUX_n9), .A2(OutputRegIn[24]), .A3(Red_done[0]), .A4(done), .ZN(Output[24]) );
  AND4_X1 Output_MUX_AND3_inst_25_U1 ( .A1(Output_MUX_n9), .A2(OutputRegIn[25]), .A3(Output_MUX_n8), .A4(Output_MUX_n10), .ZN(Output[25]) );
  AND4_X1 Output_MUX_AND3_inst_26_U1 ( .A1(Output_MUX_n9), .A2(OutputRegIn[26]), .A3(Red_done[0]), .A4(Output_MUX_n10), .ZN(Output[26]) );
  AND4_X1 Output_MUX_AND3_inst_27_U1 ( .A1(Output_MUX_n9), .A2(OutputRegIn[27]), .A3(Red_done[0]), .A4(Output_MUX_n10), .ZN(Output[27]) );
  AND4_X1 Output_MUX_AND3_inst_28_U1 ( .A1(Output_MUX_n9), .A2(OutputRegIn[28]), .A3(Output_MUX_n8), .A4(Output_MUX_n10), .ZN(Output[28]) );
  AND4_X1 Output_MUX_AND3_inst_29_U1 ( .A1(Output_MUX_n9), .A2(OutputRegIn[29]), .A3(Output_MUX_n8), .A4(Output_MUX_n10), .ZN(Output[29]) );
  AND4_X1 Output_MUX_AND3_inst_30_U1 ( .A1(Output_MUX_n9), .A2(OutputRegIn[30]), .A3(Red_done[0]), .A4(Output_MUX_n10), .ZN(Output[30]) );
  AND4_X1 Output_MUX_AND3_inst_31_U1 ( .A1(Output_MUX_n9), .A2(OutputRegIn[31]), .A3(Output_MUX_n8), .A4(Output_MUX_n10), .ZN(Output[31]) );
  AND4_X1 Output_MUX_AND3_inst_32_U1 ( .A1(Output_MUX_n9), .A2(OutputRegIn[32]), .A3(Red_done[0]), .A4(Output_MUX_n10), .ZN(Output[32]) );
  AND4_X1 Output_MUX_AND3_inst_33_U1 ( .A1(Output_MUX_n9), .A2(OutputRegIn[33]), .A3(Output_MUX_n8), .A4(Output_MUX_n10), .ZN(Output[33]) );
  AND4_X1 Output_MUX_AND3_inst_34_U1 ( .A1(Output_MUX_n9), .A2(OutputRegIn[34]), .A3(Output_MUX_n8), .A4(Output_MUX_n10), .ZN(Output[34]) );
  AND4_X1 Output_MUX_AND3_inst_35_U1 ( .A1(Output_MUX_n9), .A2(OutputRegIn[35]), .A3(Output_MUX_n8), .A4(Output_MUX_n10), .ZN(Output[35]) );
  AND4_X1 Output_MUX_AND3_inst_36_U1 ( .A1(Output_MUX_n9), .A2(OutputRegIn[36]), .A3(Output_MUX_n8), .A4(Output_MUX_n10), .ZN(Output[36]) );
  AND4_X1 Output_MUX_AND3_inst_37_U1 ( .A1(Output_MUX_n9), .A2(OutputRegIn[37]), .A3(Output_MUX_n7), .A4(done), .ZN(Output[37]) );
  AND4_X1 Output_MUX_AND3_inst_38_U1 ( .A1(Red_done[1]), .A2(OutputRegIn[38]), 
        .A3(Output_MUX_n8), .A4(done), .ZN(Output[38]) );
  AND4_X1 Output_MUX_AND3_inst_39_U1 ( .A1(Output_MUX_n9), .A2(OutputRegIn[39]), .A3(Output_MUX_n7), .A4(Output_MUX_n10), .ZN(Output[39]) );
  AND4_X1 Output_MUX_AND3_inst_40_U1 ( .A1(Output_MUX_n9), .A2(OutputRegIn[40]), .A3(Output_MUX_n8), .A4(done), .ZN(Output[40]) );
  AND4_X1 Output_MUX_AND3_inst_41_U1 ( .A1(Red_done[1]), .A2(OutputRegIn[41]), 
        .A3(Output_MUX_n7), .A4(done), .ZN(Output[41]) );
  AND4_X1 Output_MUX_AND3_inst_42_U1 ( .A1(Output_MUX_n9), .A2(OutputRegIn[42]), .A3(Output_MUX_n8), .A4(done), .ZN(Output[42]) );
  AND4_X1 Output_MUX_AND3_inst_43_U1 ( .A1(Output_MUX_n9), .A2(OutputRegIn[43]), .A3(Output_MUX_n7), .A4(Output_MUX_n10), .ZN(Output[43]) );
  AND4_X1 Output_MUX_AND3_inst_44_U1 ( .A1(Red_done[1]), .A2(OutputRegIn[44]), 
        .A3(Output_MUX_n8), .A4(done), .ZN(Output[44]) );
  AND4_X1 Output_MUX_AND3_inst_45_U1 ( .A1(Output_MUX_n9), .A2(OutputRegIn[45]), .A3(Output_MUX_n7), .A4(done), .ZN(Output[45]) );
  AND4_X1 Output_MUX_AND3_inst_46_U1 ( .A1(Output_MUX_n9), .A2(OutputRegIn[46]), .A3(Output_MUX_n8), .A4(Output_MUX_n10), .ZN(Output[46]) );
  AND4_X1 Output_MUX_AND3_inst_47_U1 ( .A1(Output_MUX_n9), .A2(OutputRegIn[47]), .A3(Output_MUX_n7), .A4(Output_MUX_n10), .ZN(Output[47]) );
  AND4_X1 Output_MUX_AND3_inst_48_U1 ( .A1(Output_MUX_n9), .A2(OutputRegIn[48]), .A3(Output_MUX_n8), .A4(done), .ZN(Output[48]) );
  AND4_X1 Output_MUX_AND3_inst_49_U1 ( .A1(Red_done[1]), .A2(OutputRegIn[49]), 
        .A3(Output_MUX_n7), .A4(done), .ZN(Output[49]) );
  AND4_X1 Output_MUX_AND3_inst_50_U1 ( .A1(Output_MUX_n9), .A2(OutputRegIn[50]), .A3(Output_MUX_n7), .A4(done), .ZN(Output[50]) );
  AND4_X1 Output_MUX_AND3_inst_51_U1 ( .A1(Output_MUX_n9), .A2(OutputRegIn[51]), .A3(Output_MUX_n7), .A4(Output_MUX_n10), .ZN(Output[51]) );
  AND4_X1 Output_MUX_AND3_inst_52_U1 ( .A1(Red_done[1]), .A2(OutputRegIn[52]), 
        .A3(Output_MUX_n7), .A4(done), .ZN(Output[52]) );
  AND4_X1 Output_MUX_AND3_inst_53_U1 ( .A1(Output_MUX_n9), .A2(OutputRegIn[53]), .A3(Output_MUX_n7), .A4(done), .ZN(Output[53]) );
  AND4_X1 Output_MUX_AND3_inst_54_U1 ( .A1(Output_MUX_n9), .A2(OutputRegIn[54]), .A3(Output_MUX_n7), .A4(Output_MUX_n10), .ZN(Output[54]) );
  AND4_X1 Output_MUX_AND3_inst_55_U1 ( .A1(Red_done[1]), .A2(OutputRegIn[55]), 
        .A3(Output_MUX_n7), .A4(done), .ZN(Output[55]) );
  AND4_X1 Output_MUX_AND3_inst_56_U1 ( .A1(Output_MUX_n9), .A2(OutputRegIn[56]), .A3(Output_MUX_n7), .A4(done), .ZN(Output[56]) );
  AND4_X1 Output_MUX_AND3_inst_57_U1 ( .A1(Output_MUX_n9), .A2(OutputRegIn[57]), .A3(Output_MUX_n7), .A4(Output_MUX_n10), .ZN(Output[57]) );
  AND4_X1 Output_MUX_AND3_inst_58_U1 ( .A1(Red_done[1]), .A2(OutputRegIn[58]), 
        .A3(Output_MUX_n7), .A4(done), .ZN(Output[58]) );
  AND4_X1 Output_MUX_AND3_inst_59_U1 ( .A1(Output_MUX_n9), .A2(OutputRegIn[59]), .A3(Output_MUX_n7), .A4(done), .ZN(Output[59]) );
  AND4_X1 Output_MUX_AND3_inst_60_U1 ( .A1(Red_done[1]), .A2(OutputRegIn[60]), 
        .A3(Output_MUX_n7), .A4(Output_MUX_n10), .ZN(Output[60]) );
  AND4_X1 Output_MUX_AND3_inst_61_U1 ( .A1(Output_MUX_n9), .A2(OutputRegIn[61]), .A3(Output_MUX_n8), .A4(done), .ZN(Output[61]) );
  AND4_X1 Output_MUX_AND3_inst_62_U1 ( .A1(Output_MUX_n9), .A2(OutputRegIn[62]), .A3(Output_MUX_n8), .A4(done), .ZN(Output[62]) );
  AND4_X1 Output_MUX_AND3_inst_63_U1 ( .A1(Output_MUX_n9), .A2(OutputRegIn[63]), .A3(Output_MUX_n8), .A4(done), .ZN(Output[63]) );
endmodule

